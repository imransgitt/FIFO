module fifo ( gnd, vdd, clk, reset, d_in, wr_en, rd_en, full, empty, d_out, fifo_counter);

input gnd, vdd;
input clk;
input reset;
input wr_en;
input rd_en;
output full;
output empty;
input [7:0] d_in;
output [7:0] d_out;
output [4:0] fifo_counter;

BUFX4 BUFX4_1 ( .gnd(gnd), .vdd(vdd), .A(_156_), .Y(_156__bF_buf5) );
BUFX4 BUFX4_2 ( .gnd(gnd), .vdd(vdd), .A(_156_), .Y(_156__bF_buf4) );
BUFX4 BUFX4_3 ( .gnd(gnd), .vdd(vdd), .A(_156_), .Y(_156__bF_buf3) );
BUFX4 BUFX4_4 ( .gnd(gnd), .vdd(vdd), .A(_156_), .Y(_156__bF_buf2) );
BUFX4 BUFX4_5 ( .gnd(gnd), .vdd(vdd), .A(_156_), .Y(_156__bF_buf1) );
BUFX4 BUFX4_6 ( .gnd(gnd), .vdd(vdd), .A(_156_), .Y(_156__bF_buf0) );
CLKBUF1 CLKBUF1_1 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf11) );
CLKBUF1 CLKBUF1_2 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf10) );
CLKBUF1 CLKBUF1_3 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf9) );
CLKBUF1 CLKBUF1_4 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf8) );
CLKBUF1 CLKBUF1_5 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf7) );
CLKBUF1 CLKBUF1_6 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf6) );
CLKBUF1 CLKBUF1_7 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf5) );
CLKBUF1 CLKBUF1_8 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf4) );
CLKBUF1 CLKBUF1_9 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf3) );
CLKBUF1 CLKBUF1_10 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf2) );
CLKBUF1 CLKBUF1_11 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf1) );
CLKBUF1 CLKBUF1_12 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf0) );
BUFX4 BUFX4_7 ( .gnd(gnd), .vdd(vdd), .A(_141_), .Y(_141__bF_buf4) );
BUFX4 BUFX4_8 ( .gnd(gnd), .vdd(vdd), .A(_141_), .Y(_141__bF_buf3) );
BUFX4 BUFX4_9 ( .gnd(gnd), .vdd(vdd), .A(_141_), .Y(_141__bF_buf2) );
BUFX4 BUFX4_10 ( .gnd(gnd), .vdd(vdd), .A(_141_), .Y(_141__bF_buf1) );
BUFX4 BUFX4_11 ( .gnd(gnd), .vdd(vdd), .A(_141_), .Y(_141__bF_buf0) );
BUFX4 BUFX4_12 ( .gnd(gnd), .vdd(vdd), .A(_132_), .Y(_132__bF_buf3) );
BUFX4 BUFX4_13 ( .gnd(gnd), .vdd(vdd), .A(_132_), .Y(_132__bF_buf2) );
BUFX4 BUFX4_14 ( .gnd(gnd), .vdd(vdd), .A(_132_), .Y(_132__bF_buf1) );
BUFX4 BUFX4_15 ( .gnd(gnd), .vdd(vdd), .A(_132_), .Y(_132__bF_buf0) );
BUFX4 BUFX4_16 ( .gnd(gnd), .vdd(vdd), .A(rd_ptr_1_), .Y(rd_ptr_1_bF_buf3_) );
BUFX4 BUFX4_17 ( .gnd(gnd), .vdd(vdd), .A(rd_ptr_1_), .Y(rd_ptr_1_bF_buf2_) );
BUFX4 BUFX4_18 ( .gnd(gnd), .vdd(vdd), .A(rd_ptr_1_), .Y(rd_ptr_1_bF_buf1_) );
BUFX4 BUFX4_19 ( .gnd(gnd), .vdd(vdd), .A(rd_ptr_1_), .Y(rd_ptr_1_bF_buf0_) );
BUFX4 BUFX4_20 ( .gnd(gnd), .vdd(vdd), .A(_155_), .Y(_155__bF_buf5) );
BUFX4 BUFX4_21 ( .gnd(gnd), .vdd(vdd), .A(_155_), .Y(_155__bF_buf4) );
BUFX4 BUFX4_22 ( .gnd(gnd), .vdd(vdd), .A(_155_), .Y(_155__bF_buf3) );
BUFX4 BUFX4_23 ( .gnd(gnd), .vdd(vdd), .A(_155_), .Y(_155__bF_buf2) );
BUFX4 BUFX4_24 ( .gnd(gnd), .vdd(vdd), .A(_155_), .Y(_155__bF_buf1) );
BUFX4 BUFX4_25 ( .gnd(gnd), .vdd(vdd), .A(_155_), .Y(_155__bF_buf0) );
BUFX4 BUFX4_26 ( .gnd(gnd), .vdd(vdd), .A(_160_), .Y(_160__bF_buf7) );
BUFX4 BUFX4_27 ( .gnd(gnd), .vdd(vdd), .A(_160_), .Y(_160__bF_buf6) );
BUFX4 BUFX4_28 ( .gnd(gnd), .vdd(vdd), .A(_160_), .Y(_160__bF_buf5) );
BUFX4 BUFX4_29 ( .gnd(gnd), .vdd(vdd), .A(_160_), .Y(_160__bF_buf4) );
BUFX4 BUFX4_30 ( .gnd(gnd), .vdd(vdd), .A(_160_), .Y(_160__bF_buf3) );
BUFX4 BUFX4_31 ( .gnd(gnd), .vdd(vdd), .A(_160_), .Y(_160__bF_buf2) );
BUFX4 BUFX4_32 ( .gnd(gnd), .vdd(vdd), .A(_160_), .Y(_160__bF_buf1) );
BUFX4 BUFX4_33 ( .gnd(gnd), .vdd(vdd), .A(_160_), .Y(_160__bF_buf0) );
BUFX4 BUFX4_34 ( .gnd(gnd), .vdd(vdd), .A(rd_ptr_3_), .Y(rd_ptr_3_bF_buf3_) );
BUFX4 BUFX4_35 ( .gnd(gnd), .vdd(vdd), .A(rd_ptr_3_), .Y(rd_ptr_3_bF_buf2_) );
BUFX4 BUFX4_36 ( .gnd(gnd), .vdd(vdd), .A(rd_ptr_3_), .Y(rd_ptr_3_bF_buf1_) );
BUFX4 BUFX4_37 ( .gnd(gnd), .vdd(vdd), .A(rd_ptr_3_), .Y(rd_ptr_3_bF_buf0_) );
BUFX4 BUFX4_38 ( .gnd(gnd), .vdd(vdd), .A(rd_ptr_0_), .Y(rd_ptr_0_bF_buf5_) );
BUFX4 BUFX4_39 ( .gnd(gnd), .vdd(vdd), .A(rd_ptr_0_), .Y(rd_ptr_0_bF_buf4_) );
BUFX4 BUFX4_40 ( .gnd(gnd), .vdd(vdd), .A(rd_ptr_0_), .Y(rd_ptr_0_bF_buf3_) );
BUFX4 BUFX4_41 ( .gnd(gnd), .vdd(vdd), .A(rd_ptr_0_), .Y(rd_ptr_0_bF_buf2_) );
BUFX4 BUFX4_42 ( .gnd(gnd), .vdd(vdd), .A(rd_ptr_0_), .Y(rd_ptr_0_bF_buf1_) );
BUFX4 BUFX4_43 ( .gnd(gnd), .vdd(vdd), .A(rd_ptr_0_), .Y(rd_ptr_0_bF_buf0_) );
BUFX4 BUFX4_44 ( .gnd(gnd), .vdd(vdd), .A(_171_), .Y(_171__bF_buf3) );
BUFX4 BUFX4_45 ( .gnd(gnd), .vdd(vdd), .A(_171_), .Y(_171__bF_buf2) );
BUFX4 BUFX4_46 ( .gnd(gnd), .vdd(vdd), .A(_171_), .Y(_171__bF_buf1) );
BUFX4 BUFX4_47 ( .gnd(gnd), .vdd(vdd), .A(_171_), .Y(_171__bF_buf0) );
MUX2X1 MUX2X1_1 ( .gnd(gnd), .vdd(vdd), .A(_455_), .B(_204_), .S(_488_), .Y(_100_) );
MUX2X1 MUX2X1_2 ( .gnd(gnd), .vdd(vdd), .A(_459_), .B(_234_), .S(_488_), .Y(_101_) );
NOR2X1 NOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(memory_6__2_), .B(_488_), .Y(_489_) );
AOI21X1 AOI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(_461_), .B(_488_), .C(_489_), .Y(_102_) );
MUX2X1 MUX2X1_3 ( .gnd(gnd), .vdd(vdd), .A(_463_), .B(_288_), .S(_488_), .Y(_103_) );
MUX2X1 MUX2X1_4 ( .gnd(gnd), .vdd(vdd), .A(_465_), .B(_316_), .S(_488_), .Y(_104_) );
MUX2X1 MUX2X1_5 ( .gnd(gnd), .vdd(vdd), .A(_467_), .B(_344_), .S(_488_), .Y(_105_) );
MUX2X1 MUX2X1_6 ( .gnd(gnd), .vdd(vdd), .A(_469_), .B(_372_), .S(_488_), .Y(_106_) );
MUX2X1 MUX2X1_7 ( .gnd(gnd), .vdd(vdd), .A(_471_), .B(_400_), .S(_488_), .Y(_107_) );
NAND2X1 NAND2X1_1 ( .gnd(gnd), .vdd(vdd), .A(memory_7__0_), .B(_171__bF_buf3), .Y(_490_) );
OAI21X1 OAI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(_171__bF_buf2), .B(_431_), .C(_490_), .Y(_108_) );
NAND2X1 NAND2X1_2 ( .gnd(gnd), .vdd(vdd), .A(memory_7__1_), .B(_171__bF_buf1), .Y(_491_) );
OAI21X1 OAI21X1_2 ( .gnd(gnd), .vdd(vdd), .A(_171__bF_buf0), .B(_433_), .C(_491_), .Y(_109_) );
NAND2X1 NAND2X1_3 ( .gnd(gnd), .vdd(vdd), .A(memory_7__2_), .B(_171__bF_buf3), .Y(_492_) );
OAI21X1 OAI21X1_3 ( .gnd(gnd), .vdd(vdd), .A(_171__bF_buf2), .B(_435_), .C(_492_), .Y(_110_) );
NAND2X1 NAND2X1_4 ( .gnd(gnd), .vdd(vdd), .A(memory_7__3_), .B(_171__bF_buf1), .Y(_493_) );
OAI21X1 OAI21X1_4 ( .gnd(gnd), .vdd(vdd), .A(_171__bF_buf0), .B(_437_), .C(_493_), .Y(_111_) );
NAND2X1 NAND2X1_5 ( .gnd(gnd), .vdd(vdd), .A(memory_7__4_), .B(_171__bF_buf3), .Y(_494_) );
OAI21X1 OAI21X1_5 ( .gnd(gnd), .vdd(vdd), .A(_171__bF_buf2), .B(_439_), .C(_494_), .Y(_112_) );
NAND2X1 NAND2X1_6 ( .gnd(gnd), .vdd(vdd), .A(memory_7__5_), .B(_171__bF_buf1), .Y(_495_) );
OAI21X1 OAI21X1_6 ( .gnd(gnd), .vdd(vdd), .A(_171__bF_buf0), .B(_441_), .C(_495_), .Y(_113_) );
NAND2X1 NAND2X1_7 ( .gnd(gnd), .vdd(vdd), .A(memory_7__6_), .B(_171__bF_buf3), .Y(_496_) );
OAI21X1 OAI21X1_7 ( .gnd(gnd), .vdd(vdd), .A(_171__bF_buf2), .B(_443_), .C(_496_), .Y(_114_) );
NAND2X1 NAND2X1_8 ( .gnd(gnd), .vdd(vdd), .A(memory_7__7_), .B(_171__bF_buf1), .Y(_497_) );
OAI21X1 OAI21X1_8 ( .gnd(gnd), .vdd(vdd), .A(_146_), .B(_171__bF_buf0), .C(_497_), .Y(_115_) );
NOR2X1 NOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(wr_ptr_2_), .B(_138_), .Y(_498_) );
NAND2X1 NAND2X1_9 ( .gnd(gnd), .vdd(vdd), .A(_429_), .B(_498_), .Y(_499_) );
NOR2X1 NOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(_499_), .B(_149_), .Y(_500_) );
NOR2X1 NOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(memory_8__0_), .B(_500_), .Y(_501_) );
AOI21X1 AOI21X1_2 ( .gnd(gnd), .vdd(vdd), .A(_455_), .B(_500_), .C(_501_), .Y(_116_) );
NOR2X1 NOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(memory_8__1_), .B(_500_), .Y(_502_) );
AOI21X1 AOI21X1_3 ( .gnd(gnd), .vdd(vdd), .A(_459_), .B(_500_), .C(_502_), .Y(_117_) );
NOR2X1 NOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(memory_8__2_), .B(_500_), .Y(_503_) );
AOI21X1 AOI21X1_4 ( .gnd(gnd), .vdd(vdd), .A(_461_), .B(_500_), .C(_503_), .Y(_118_) );
NOR2X1 NOR2X1_7 ( .gnd(gnd), .vdd(vdd), .A(memory_8__3_), .B(_500_), .Y(_504_) );
AOI21X1 AOI21X1_5 ( .gnd(gnd), .vdd(vdd), .A(_463_), .B(_500_), .C(_504_), .Y(_119_) );
NOR2X1 NOR2X1_8 ( .gnd(gnd), .vdd(vdd), .A(memory_8__4_), .B(_500_), .Y(_505_) );
AOI21X1 AOI21X1_6 ( .gnd(gnd), .vdd(vdd), .A(_465_), .B(_500_), .C(_505_), .Y(_120_) );
NOR2X1 NOR2X1_9 ( .gnd(gnd), .vdd(vdd), .A(memory_8__5_), .B(_500_), .Y(_506_) );
AOI21X1 AOI21X1_7 ( .gnd(gnd), .vdd(vdd), .A(_467_), .B(_500_), .C(_506_), .Y(_121_) );
NOR2X1 NOR2X1_10 ( .gnd(gnd), .vdd(vdd), .A(memory_8__6_), .B(_500_), .Y(_507_) );
AOI21X1 AOI21X1_8 ( .gnd(gnd), .vdd(vdd), .A(_469_), .B(_500_), .C(_507_), .Y(_122_) );
NOR2X1 NOR2X1_11 ( .gnd(gnd), .vdd(vdd), .A(memory_8__7_), .B(_500_), .Y(_508_) );
AOI21X1 AOI21X1_9 ( .gnd(gnd), .vdd(vdd), .A(_471_), .B(_500_), .C(_508_), .Y(_123_) );
NAND2X1 NAND2X1_10 ( .gnd(gnd), .vdd(vdd), .A(_167_), .B(_498_), .Y(_509_) );
NOR2X1 NOR2X1_12 ( .gnd(gnd), .vdd(vdd), .A(_509_), .B(_149_), .Y(_510_) );
NOR2X1 NOR2X1_13 ( .gnd(gnd), .vdd(vdd), .A(memory_9__0_), .B(_510_), .Y(_511_) );
AOI21X1 AOI21X1_10 ( .gnd(gnd), .vdd(vdd), .A(_431_), .B(_510_), .C(_511_), .Y(_124_) );
NOR2X1 NOR2X1_14 ( .gnd(gnd), .vdd(vdd), .A(memory_9__1_), .B(_510_), .Y(_512_) );
AOI21X1 AOI21X1_11 ( .gnd(gnd), .vdd(vdd), .A(_433_), .B(_510_), .C(_512_), .Y(_125_) );
NOR2X1 NOR2X1_15 ( .gnd(gnd), .vdd(vdd), .A(memory_9__2_), .B(_510_), .Y(_513_) );
AOI21X1 AOI21X1_12 ( .gnd(gnd), .vdd(vdd), .A(_435_), .B(_510_), .C(_513_), .Y(_126_) );
NOR2X1 NOR2X1_16 ( .gnd(gnd), .vdd(vdd), .A(memory_9__3_), .B(_510_), .Y(_514_) );
AOI21X1 AOI21X1_13 ( .gnd(gnd), .vdd(vdd), .A(_437_), .B(_510_), .C(_514_), .Y(_127_) );
NOR2X1 NOR2X1_17 ( .gnd(gnd), .vdd(vdd), .A(memory_9__4_), .B(_510_), .Y(_515_) );
AOI21X1 AOI21X1_14 ( .gnd(gnd), .vdd(vdd), .A(_439_), .B(_510_), .C(_515_), .Y(_128_) );
NOR2X1 NOR2X1_18 ( .gnd(gnd), .vdd(vdd), .A(memory_9__5_), .B(_510_), .Y(_516_) );
AOI21X1 AOI21X1_15 ( .gnd(gnd), .vdd(vdd), .A(_441_), .B(_510_), .C(_516_), .Y(_129_) );
NOR2X1 NOR2X1_19 ( .gnd(gnd), .vdd(vdd), .A(memory_9__6_), .B(_510_), .Y(_517_) );
AOI21X1 AOI21X1_16 ( .gnd(gnd), .vdd(vdd), .A(_443_), .B(_510_), .C(_517_), .Y(_130_) );
NOR2X1 NOR2X1_20 ( .gnd(gnd), .vdd(vdd), .A(memory_9__7_), .B(_510_), .Y(_518_) );
AOI21X1 AOI21X1_17 ( .gnd(gnd), .vdd(vdd), .A(_146_), .B(_510_), .C(_518_), .Y(_131_) );
NAND2X1 NAND2X1_11 ( .gnd(gnd), .vdd(vdd), .A(_166_), .B(_498_), .Y(_519_) );
NOR2X1 NOR2X1_21 ( .gnd(gnd), .vdd(vdd), .A(_519_), .B(_149_), .Y(_520_) );
MUX2X1 MUX2X1_8 ( .gnd(gnd), .vdd(vdd), .A(_455_), .B(_226_), .S(_520_), .Y(_12_) );
NOR2X1 NOR2X1_22 ( .gnd(gnd), .vdd(vdd), .A(memory_10__1_), .B(_520_), .Y(_521_) );
AOI21X1 AOI21X1_18 ( .gnd(gnd), .vdd(vdd), .A(_459_), .B(_520_), .C(_521_), .Y(_13_) );
NOR2X1 NOR2X1_23 ( .gnd(gnd), .vdd(vdd), .A(memory_10__2_), .B(_520_), .Y(_522_) );
AOI21X1 AOI21X1_19 ( .gnd(gnd), .vdd(vdd), .A(_461_), .B(_520_), .C(_522_), .Y(_14_) );
MUX2X1 MUX2X1_9 ( .gnd(gnd), .vdd(vdd), .A(_463_), .B(_303_), .S(_520_), .Y(_15_) );
MUX2X1 MUX2X1_10 ( .gnd(gnd), .vdd(vdd), .A(_465_), .B(_331_), .S(_520_), .Y(_16_) );
NOR2X1 NOR2X1_24 ( .gnd(gnd), .vdd(vdd), .A(memory_10__5_), .B(_520_), .Y(_523_) );
AOI21X1 AOI21X1_20 ( .gnd(gnd), .vdd(vdd), .A(_467_), .B(_520_), .C(_523_), .Y(_17_) );
MUX2X1 MUX2X1_11 ( .gnd(gnd), .vdd(vdd), .A(_469_), .B(_387_), .S(_520_), .Y(_18_) );
NOR2X1 NOR2X1_25 ( .gnd(gnd), .vdd(vdd), .A(memory_10__7_), .B(_520_), .Y(_524_) );
AOI21X1 AOI21X1_21 ( .gnd(gnd), .vdd(vdd), .A(_471_), .B(_520_), .C(_524_), .Y(_19_) );
NAND3X1 NAND3X1_1 ( .gnd(gnd), .vdd(vdd), .A(_144_), .B(_498_), .C(_141__bF_buf4), .Y(_525_) );
NAND2X1 NAND2X1_12 ( .gnd(gnd), .vdd(vdd), .A(memory_11__0_), .B(_525_), .Y(_526_) );
OAI21X1 OAI21X1_9 ( .gnd(gnd), .vdd(vdd), .A(_431_), .B(_525_), .C(_526_), .Y(_20_) );
NAND2X1 NAND2X1_13 ( .gnd(gnd), .vdd(vdd), .A(memory_11__1_), .B(_525_), .Y(_527_) );
OAI21X1 OAI21X1_10 ( .gnd(gnd), .vdd(vdd), .A(_433_), .B(_525_), .C(_527_), .Y(_21_) );
NAND2X1 NAND2X1_14 ( .gnd(gnd), .vdd(vdd), .A(memory_11__2_), .B(_525_), .Y(_528_) );
OAI21X1 OAI21X1_11 ( .gnd(gnd), .vdd(vdd), .A(_435_), .B(_525_), .C(_528_), .Y(_22_) );
NAND2X1 NAND2X1_15 ( .gnd(gnd), .vdd(vdd), .A(memory_11__3_), .B(_525_), .Y(_529_) );
OAI21X1 OAI21X1_12 ( .gnd(gnd), .vdd(vdd), .A(_437_), .B(_525_), .C(_529_), .Y(_23_) );
NAND2X1 NAND2X1_16 ( .gnd(gnd), .vdd(vdd), .A(memory_11__4_), .B(_525_), .Y(_530_) );
OAI21X1 OAI21X1_13 ( .gnd(gnd), .vdd(vdd), .A(_439_), .B(_525_), .C(_530_), .Y(_24_) );
NAND2X1 NAND2X1_17 ( .gnd(gnd), .vdd(vdd), .A(memory_11__5_), .B(_525_), .Y(_531_) );
OAI21X1 OAI21X1_14 ( .gnd(gnd), .vdd(vdd), .A(_441_), .B(_525_), .C(_531_), .Y(_25_) );
NAND2X1 NAND2X1_18 ( .gnd(gnd), .vdd(vdd), .A(memory_11__6_), .B(_525_), .Y(_532_) );
OAI21X1 OAI21X1_15 ( .gnd(gnd), .vdd(vdd), .A(_443_), .B(_525_), .C(_532_), .Y(_26_) );
NAND2X1 NAND2X1_19 ( .gnd(gnd), .vdd(vdd), .A(memory_11__7_), .B(_525_), .Y(_533_) );
OAI21X1 OAI21X1_16 ( .gnd(gnd), .vdd(vdd), .A(_146_), .B(_525_), .C(_533_), .Y(_27_) );
NAND3X1 NAND3X1_2 ( .gnd(gnd), .vdd(vdd), .A(_140_), .B(_429_), .C(_141__bF_buf3), .Y(_534_) );
NAND2X1 NAND2X1_20 ( .gnd(gnd), .vdd(vdd), .A(memory_12__0_), .B(_534_), .Y(_535_) );
OAI21X1 OAI21X1_17 ( .gnd(gnd), .vdd(vdd), .A(_431_), .B(_534_), .C(_535_), .Y(_28_) );
NAND2X1 NAND2X1_21 ( .gnd(gnd), .vdd(vdd), .A(memory_12__1_), .B(_534_), .Y(_536_) );
OAI21X1 OAI21X1_18 ( .gnd(gnd), .vdd(vdd), .A(_433_), .B(_534_), .C(_536_), .Y(_29_) );
NAND2X1 NAND2X1_22 ( .gnd(gnd), .vdd(vdd), .A(memory_12__2_), .B(_534_), .Y(_537_) );
OAI21X1 OAI21X1_19 ( .gnd(gnd), .vdd(vdd), .A(_435_), .B(_534_), .C(_537_), .Y(_30_) );
NAND2X1 NAND2X1_23 ( .gnd(gnd), .vdd(vdd), .A(memory_12__3_), .B(_534_), .Y(_538_) );
OAI21X1 OAI21X1_20 ( .gnd(gnd), .vdd(vdd), .A(_437_), .B(_534_), .C(_538_), .Y(_31_) );
NAND2X1 NAND2X1_24 ( .gnd(gnd), .vdd(vdd), .A(memory_12__4_), .B(_534_), .Y(_539_) );
OAI21X1 OAI21X1_21 ( .gnd(gnd), .vdd(vdd), .A(_439_), .B(_534_), .C(_539_), .Y(_32_) );
NAND2X1 NAND2X1_25 ( .gnd(gnd), .vdd(vdd), .A(memory_12__5_), .B(_534_), .Y(_540_) );
OAI21X1 OAI21X1_22 ( .gnd(gnd), .vdd(vdd), .A(_441_), .B(_534_), .C(_540_), .Y(_33_) );
NAND2X1 NAND2X1_26 ( .gnd(gnd), .vdd(vdd), .A(memory_12__6_), .B(_534_), .Y(_541_) );
OAI21X1 OAI21X1_23 ( .gnd(gnd), .vdd(vdd), .A(_443_), .B(_534_), .C(_541_), .Y(_34_) );
NAND2X1 NAND2X1_27 ( .gnd(gnd), .vdd(vdd), .A(memory_12__7_), .B(_534_), .Y(_542_) );
OAI21X1 OAI21X1_24 ( .gnd(gnd), .vdd(vdd), .A(_146_), .B(_534_), .C(_542_), .Y(_35_) );
NAND3X1 NAND3X1_3 ( .gnd(gnd), .vdd(vdd), .A(_140_), .B(_167_), .C(_141__bF_buf2), .Y(_543_) );
NAND2X1 NAND2X1_28 ( .gnd(gnd), .vdd(vdd), .A(memory_13__0_), .B(_543_), .Y(_544_) );
OAI21X1 OAI21X1_25 ( .gnd(gnd), .vdd(vdd), .A(_431_), .B(_543_), .C(_544_), .Y(_36_) );
NAND2X1 NAND2X1_29 ( .gnd(gnd), .vdd(vdd), .A(memory_13__1_), .B(_543_), .Y(_545_) );
OAI21X1 OAI21X1_26 ( .gnd(gnd), .vdd(vdd), .A(_433_), .B(_543_), .C(_545_), .Y(_37_) );
NAND2X1 NAND2X1_30 ( .gnd(gnd), .vdd(vdd), .A(memory_13__2_), .B(_543_), .Y(_546_) );
OAI21X1 OAI21X1_27 ( .gnd(gnd), .vdd(vdd), .A(_435_), .B(_543_), .C(_546_), .Y(_38_) );
NAND2X1 NAND2X1_31 ( .gnd(gnd), .vdd(vdd), .A(memory_13__3_), .B(_543_), .Y(_547_) );
OAI21X1 OAI21X1_28 ( .gnd(gnd), .vdd(vdd), .A(_437_), .B(_543_), .C(_547_), .Y(_39_) );
NAND2X1 NAND2X1_32 ( .gnd(gnd), .vdd(vdd), .A(memory_13__4_), .B(_543_), .Y(_548_) );
OAI21X1 OAI21X1_29 ( .gnd(gnd), .vdd(vdd), .A(_439_), .B(_543_), .C(_548_), .Y(_40_) );
NAND2X1 NAND2X1_33 ( .gnd(gnd), .vdd(vdd), .A(memory_13__5_), .B(_543_), .Y(_549_) );
OAI21X1 OAI21X1_30 ( .gnd(gnd), .vdd(vdd), .A(_441_), .B(_543_), .C(_549_), .Y(_41_) );
NAND2X1 NAND2X1_34 ( .gnd(gnd), .vdd(vdd), .A(memory_13__6_), .B(_543_), .Y(_550_) );
OAI21X1 OAI21X1_31 ( .gnd(gnd), .vdd(vdd), .A(_443_), .B(_543_), .C(_550_), .Y(_42_) );
NAND2X1 NAND2X1_35 ( .gnd(gnd), .vdd(vdd), .A(memory_13__7_), .B(_543_), .Y(_551_) );
OAI21X1 OAI21X1_32 ( .gnd(gnd), .vdd(vdd), .A(_146_), .B(_543_), .C(_551_), .Y(_43_) );
NAND3X1 NAND3X1_4 ( .gnd(gnd), .vdd(vdd), .A(_140_), .B(_166_), .C(_141__bF_buf1), .Y(_552_) );
NAND2X1 NAND2X1_36 ( .gnd(gnd), .vdd(vdd), .A(memory_14__0_), .B(_552_), .Y(_553_) );
OAI21X1 OAI21X1_33 ( .gnd(gnd), .vdd(vdd), .A(_431_), .B(_552_), .C(_553_), .Y(_44_) );
NAND2X1 NAND2X1_37 ( .gnd(gnd), .vdd(vdd), .A(memory_14__1_), .B(_552_), .Y(_554_) );
OAI21X1 OAI21X1_34 ( .gnd(gnd), .vdd(vdd), .A(_433_), .B(_552_), .C(_554_), .Y(_45_) );
NAND2X1 NAND2X1_38 ( .gnd(gnd), .vdd(vdd), .A(memory_14__2_), .B(_552_), .Y(_555_) );
OAI21X1 OAI21X1_35 ( .gnd(gnd), .vdd(vdd), .A(_435_), .B(_552_), .C(_555_), .Y(_46_) );
NAND2X1 NAND2X1_39 ( .gnd(gnd), .vdd(vdd), .A(memory_14__3_), .B(_552_), .Y(_556_) );
OAI21X1 OAI21X1_36 ( .gnd(gnd), .vdd(vdd), .A(_437_), .B(_552_), .C(_556_), .Y(_47_) );
NAND2X1 NAND2X1_40 ( .gnd(gnd), .vdd(vdd), .A(memory_14__4_), .B(_552_), .Y(_557_) );
OAI21X1 OAI21X1_37 ( .gnd(gnd), .vdd(vdd), .A(_439_), .B(_552_), .C(_557_), .Y(_48_) );
NAND2X1 NAND2X1_41 ( .gnd(gnd), .vdd(vdd), .A(memory_14__5_), .B(_552_), .Y(_558_) );
OAI21X1 OAI21X1_38 ( .gnd(gnd), .vdd(vdd), .A(_441_), .B(_552_), .C(_558_), .Y(_49_) );
NAND2X1 NAND2X1_42 ( .gnd(gnd), .vdd(vdd), .A(memory_14__6_), .B(_552_), .Y(_559_) );
OAI21X1 OAI21X1_39 ( .gnd(gnd), .vdd(vdd), .A(_443_), .B(_552_), .C(_559_), .Y(_50_) );
NAND2X1 NAND2X1_43 ( .gnd(gnd), .vdd(vdd), .A(memory_14__7_), .B(_552_), .Y(_560_) );
OAI21X1 OAI21X1_40 ( .gnd(gnd), .vdd(vdd), .A(_146_), .B(_552_), .C(_560_), .Y(_51_) );
NAND2X1 NAND2X1_44 ( .gnd(gnd), .vdd(vdd), .A(memory_15__0_), .B(_145_), .Y(_561_) );
OAI21X1 OAI21X1_41 ( .gnd(gnd), .vdd(vdd), .A(_145_), .B(_431_), .C(_561_), .Y(_52_) );
NAND2X1 NAND2X1_45 ( .gnd(gnd), .vdd(vdd), .A(memory_15__1_), .B(_145_), .Y(_562_) );
OAI21X1 OAI21X1_42 ( .gnd(gnd), .vdd(vdd), .A(_145_), .B(_433_), .C(_562_), .Y(_53_) );
NAND2X1 NAND2X1_46 ( .gnd(gnd), .vdd(vdd), .A(memory_15__2_), .B(_145_), .Y(_563_) );
OAI21X1 OAI21X1_43 ( .gnd(gnd), .vdd(vdd), .A(_145_), .B(_435_), .C(_563_), .Y(_54_) );
NAND2X1 NAND2X1_47 ( .gnd(gnd), .vdd(vdd), .A(memory_15__3_), .B(_145_), .Y(_564_) );
OAI21X1 OAI21X1_44 ( .gnd(gnd), .vdd(vdd), .A(_145_), .B(_437_), .C(_564_), .Y(_55_) );
NAND2X1 NAND2X1_48 ( .gnd(gnd), .vdd(vdd), .A(memory_15__4_), .B(_145_), .Y(_565_) );
OAI21X1 OAI21X1_45 ( .gnd(gnd), .vdd(vdd), .A(_145_), .B(_439_), .C(_565_), .Y(_56_) );
NAND2X1 NAND2X1_49 ( .gnd(gnd), .vdd(vdd), .A(memory_15__5_), .B(_145_), .Y(_566_) );
OAI21X1 OAI21X1_46 ( .gnd(gnd), .vdd(vdd), .A(_145_), .B(_441_), .C(_566_), .Y(_57_) );
NAND2X1 NAND2X1_50 ( .gnd(gnd), .vdd(vdd), .A(memory_15__6_), .B(_145_), .Y(_567_) );
OAI21X1 OAI21X1_47 ( .gnd(gnd), .vdd(vdd), .A(_145_), .B(_443_), .C(_567_), .Y(_58_) );
INVX8 INVX8_1 ( .gnd(gnd), .vdd(vdd), .A(reset), .Y(_132_) );
BUFX2 BUFX2_1 ( .gnd(gnd), .vdd(vdd), .A(_568__0_), .Y(d_out[0]) );
BUFX2 BUFX2_2 ( .gnd(gnd), .vdd(vdd), .A(_568__1_), .Y(d_out[1]) );
BUFX2 BUFX2_3 ( .gnd(gnd), .vdd(vdd), .A(_568__2_), .Y(d_out[2]) );
BUFX2 BUFX2_4 ( .gnd(gnd), .vdd(vdd), .A(_568__3_), .Y(d_out[3]) );
BUFX2 BUFX2_5 ( .gnd(gnd), .vdd(vdd), .A(_568__4_), .Y(d_out[4]) );
BUFX2 BUFX2_6 ( .gnd(gnd), .vdd(vdd), .A(_568__5_), .Y(d_out[5]) );
BUFX2 BUFX2_7 ( .gnd(gnd), .vdd(vdd), .A(_568__6_), .Y(d_out[6]) );
BUFX2 BUFX2_8 ( .gnd(gnd), .vdd(vdd), .A(_568__7_), .Y(d_out[7]) );
BUFX2 BUFX2_9 ( .gnd(gnd), .vdd(vdd), .A(_569_), .Y(empty) );
BUFX2 BUFX2_10 ( .gnd(gnd), .vdd(vdd), .A(_570__0_), .Y(fifo_counter[0]) );
BUFX2 BUFX2_11 ( .gnd(gnd), .vdd(vdd), .A(_570__1_), .Y(fifo_counter[1]) );
BUFX2 BUFX2_12 ( .gnd(gnd), .vdd(vdd), .A(_570__2_), .Y(fifo_counter[2]) );
BUFX2 BUFX2_13 ( .gnd(gnd), .vdd(vdd), .A(_570__3_), .Y(fifo_counter[3]) );
BUFX2 BUFX2_14 ( .gnd(gnd), .vdd(vdd), .A(_570__4_), .Y(fifo_counter[4]) );
BUFX2 BUFX2_15 ( .gnd(gnd), .vdd(vdd), .A(_571_), .Y(full) );
DFFPOSX1 DFFPOSX1_1 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_76_), .Q(memory_3__0_) );
DFFPOSX1 DFFPOSX1_2 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_77_), .Q(memory_3__1_) );
DFFPOSX1 DFFPOSX1_3 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_78_), .Q(memory_3__2_) );
DFFPOSX1 DFFPOSX1_4 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_79_), .Q(memory_3__3_) );
DFFPOSX1 DFFPOSX1_5 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_80_), .Q(memory_3__4_) );
DFFPOSX1 DFFPOSX1_6 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_81_), .Q(memory_3__5_) );
DFFPOSX1 DFFPOSX1_7 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_82_), .Q(memory_3__6_) );
DFFPOSX1 DFFPOSX1_8 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_83_), .Q(memory_3__7_) );
DFFPOSX1 DFFPOSX1_9 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_84_), .Q(memory_4__0_) );
DFFPOSX1 DFFPOSX1_10 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_85_), .Q(memory_4__1_) );
DFFPOSX1 DFFPOSX1_11 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_86_), .Q(memory_4__2_) );
DFFPOSX1 DFFPOSX1_12 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_87_), .Q(memory_4__3_) );
DFFPOSX1 DFFPOSX1_13 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_88_), .Q(memory_4__4_) );
DFFPOSX1 DFFPOSX1_14 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_89_), .Q(memory_4__5_) );
DFFPOSX1 DFFPOSX1_15 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_90_), .Q(memory_4__6_) );
DFFPOSX1 DFFPOSX1_16 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_91_), .Q(memory_4__7_) );
DFFPOSX1 DFFPOSX1_17 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_60_), .Q(memory_1__0_) );
DFFPOSX1 DFFPOSX1_18 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_61_), .Q(memory_1__1_) );
DFFPOSX1 DFFPOSX1_19 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_62_), .Q(memory_1__2_) );
DFFPOSX1 DFFPOSX1_20 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_63_), .Q(memory_1__3_) );
DFFPOSX1 DFFPOSX1_21 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_64_), .Q(memory_1__4_) );
DFFPOSX1 DFFPOSX1_22 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_65_), .Q(memory_1__5_) );
DFFPOSX1 DFFPOSX1_23 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_66_), .Q(memory_1__6_) );
DFFPOSX1 DFFPOSX1_24 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_67_), .Q(memory_1__7_) );
DFFPOSX1 DFFPOSX1_25 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_12_), .Q(memory_10__0_) );
DFFPOSX1 DFFPOSX1_26 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_13_), .Q(memory_10__1_) );
DFFPOSX1 DFFPOSX1_27 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_14_), .Q(memory_10__2_) );
DFFPOSX1 DFFPOSX1_28 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_15_), .Q(memory_10__3_) );
DFFPOSX1 DFFPOSX1_29 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_16_), .Q(memory_10__4_) );
DFFPOSX1 DFFPOSX1_30 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_17_), .Q(memory_10__5_) );
DFFPOSX1 DFFPOSX1_31 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_18_), .Q(memory_10__6_) );
DFFPOSX1 DFFPOSX1_32 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_19_), .Q(memory_10__7_) );
DFFPOSX1 DFFPOSX1_33 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_108_), .Q(memory_7__0_) );
DFFPOSX1 DFFPOSX1_34 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_109_), .Q(memory_7__1_) );
DFFPOSX1 DFFPOSX1_35 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_110_), .Q(memory_7__2_) );
DFFPOSX1 DFFPOSX1_36 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_111_), .Q(memory_7__3_) );
DFFPOSX1 DFFPOSX1_37 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_112_), .Q(memory_7__4_) );
DFFPOSX1 DFFPOSX1_38 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_113_), .Q(memory_7__5_) );
DFFPOSX1 DFFPOSX1_39 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_114_), .Q(memory_7__6_) );
DFFPOSX1 DFFPOSX1_40 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_115_), .Q(memory_7__7_) );
DFFPOSX1 DFFPOSX1_41 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_124_), .Q(memory_9__0_) );
DFFPOSX1 DFFPOSX1_42 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_125_), .Q(memory_9__1_) );
DFFPOSX1 DFFPOSX1_43 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_126_), .Q(memory_9__2_) );
DFFPOSX1 DFFPOSX1_44 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_127_), .Q(memory_9__3_) );
DFFPOSX1 DFFPOSX1_45 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_128_), .Q(memory_9__4_) );
DFFPOSX1 DFFPOSX1_46 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_129_), .Q(memory_9__5_) );
DFFPOSX1 DFFPOSX1_47 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_130_), .Q(memory_9__6_) );
DFFPOSX1 DFFPOSX1_48 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_131_), .Q(memory_9__7_) );
DFFPOSX1 DFFPOSX1_49 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_100_), .Q(memory_6__0_) );
DFFPOSX1 DFFPOSX1_50 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_101_), .Q(memory_6__1_) );
DFFPOSX1 DFFPOSX1_51 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_102_), .Q(memory_6__2_) );
DFFPOSX1 DFFPOSX1_52 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_103_), .Q(memory_6__3_) );
DFFPOSX1 DFFPOSX1_53 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_104_), .Q(memory_6__4_) );
DFFPOSX1 DFFPOSX1_54 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_105_), .Q(memory_6__5_) );
DFFPOSX1 DFFPOSX1_55 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_106_), .Q(memory_6__6_) );
DFFPOSX1 DFFPOSX1_56 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_107_), .Q(memory_6__7_) );
DFFPOSX1 DFFPOSX1_57 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_4_), .Q(memory_0__0_) );
DFFPOSX1 DFFPOSX1_58 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_5_), .Q(memory_0__1_) );
DFFPOSX1 DFFPOSX1_59 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_6_), .Q(memory_0__2_) );
DFFPOSX1 DFFPOSX1_60 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_7_), .Q(memory_0__3_) );
DFFPOSX1 DFFPOSX1_61 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_8_), .Q(memory_0__4_) );
DFFPOSX1 DFFPOSX1_62 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_9_), .Q(memory_0__5_) );
DFFPOSX1 DFFPOSX1_63 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_10_), .Q(memory_0__6_) );
DFFPOSX1 DFFPOSX1_64 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_11_), .Q(memory_0__7_) );
DFFPOSX1 DFFPOSX1_65 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_68_), .Q(memory_2__0_) );
DFFPOSX1 DFFPOSX1_66 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_69_), .Q(memory_2__1_) );
DFFPOSX1 DFFPOSX1_67 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_70_), .Q(memory_2__2_) );
DFFPOSX1 DFFPOSX1_68 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_71_), .Q(memory_2__3_) );
DFFPOSX1 DFFPOSX1_69 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_72_), .Q(memory_2__4_) );
DFFPOSX1 DFFPOSX1_70 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_73_), .Q(memory_2__5_) );
DFFPOSX1 DFFPOSX1_71 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_74_), .Q(memory_2__6_) );
DFFPOSX1 DFFPOSX1_72 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_75_), .Q(memory_2__7_) );
DFFPOSX1 DFFPOSX1_73 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_116_), .Q(memory_8__0_) );
DFFPOSX1 DFFPOSX1_74 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_117_), .Q(memory_8__1_) );
DFFPOSX1 DFFPOSX1_75 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_118_), .Q(memory_8__2_) );
DFFPOSX1 DFFPOSX1_76 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_119_), .Q(memory_8__3_) );
DFFPOSX1 DFFPOSX1_77 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_120_), .Q(memory_8__4_) );
DFFPOSX1 DFFPOSX1_78 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_121_), .Q(memory_8__5_) );
DFFPOSX1 DFFPOSX1_79 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_122_), .Q(memory_8__6_) );
DFFPOSX1 DFFPOSX1_80 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_123_), .Q(memory_8__7_) );
DFFPOSX1 DFFPOSX1_81 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_52_), .Q(memory_15__0_) );
DFFPOSX1 DFFPOSX1_82 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_53_), .Q(memory_15__1_) );
DFFPOSX1 DFFPOSX1_83 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_54_), .Q(memory_15__2_) );
DFFPOSX1 DFFPOSX1_84 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_55_), .Q(memory_15__3_) );
DFFPOSX1 DFFPOSX1_85 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_56_), .Q(memory_15__4_) );
DFFPOSX1 DFFPOSX1_86 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_57_), .Q(memory_15__5_) );
DFFPOSX1 DFFPOSX1_87 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_58_), .Q(memory_15__6_) );
DFFPOSX1 DFFPOSX1_88 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_59_), .Q(memory_15__7_) );
DFFPOSX1 DFFPOSX1_89 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_44_), .Q(memory_14__0_) );
DFFPOSX1 DFFPOSX1_90 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_45_), .Q(memory_14__1_) );
DFFPOSX1 DFFPOSX1_91 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_46_), .Q(memory_14__2_) );
DFFPOSX1 DFFPOSX1_92 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_47_), .Q(memory_14__3_) );
DFFPOSX1 DFFPOSX1_93 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_48_), .Q(memory_14__4_) );
DFFPOSX1 DFFPOSX1_94 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_49_), .Q(memory_14__5_) );
DFFPOSX1 DFFPOSX1_95 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_50_), .Q(memory_14__6_) );
DFFPOSX1 DFFPOSX1_96 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_51_), .Q(memory_14__7_) );
DFFPOSX1 DFFPOSX1_97 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_92_), .Q(memory_5__0_) );
DFFPOSX1 DFFPOSX1_98 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_93_), .Q(memory_5__1_) );
DFFPOSX1 DFFPOSX1_99 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_94_), .Q(memory_5__2_) );
DFFPOSX1 DFFPOSX1_100 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_95_), .Q(memory_5__3_) );
DFFPOSX1 DFFPOSX1_101 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_96_), .Q(memory_5__4_) );
DFFPOSX1 DFFPOSX1_102 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_97_), .Q(memory_5__5_) );
DFFPOSX1 DFFPOSX1_103 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_98_), .Q(memory_5__6_) );
DFFPOSX1 DFFPOSX1_104 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_99_), .Q(memory_5__7_) );
DFFPOSX1 DFFPOSX1_105 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_36_), .Q(memory_13__0_) );
DFFPOSX1 DFFPOSX1_106 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_37_), .Q(memory_13__1_) );
DFFPOSX1 DFFPOSX1_107 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_38_), .Q(memory_13__2_) );
DFFPOSX1 DFFPOSX1_108 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_39_), .Q(memory_13__3_) );
DFFPOSX1 DFFPOSX1_109 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_40_), .Q(memory_13__4_) );
DFFPOSX1 DFFPOSX1_110 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_41_), .Q(memory_13__5_) );
DFFPOSX1 DFFPOSX1_111 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_42_), .Q(memory_13__6_) );
DFFPOSX1 DFFPOSX1_112 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_43_), .Q(memory_13__7_) );
DFFPOSX1 DFFPOSX1_113 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_28_), .Q(memory_12__0_) );
DFFPOSX1 DFFPOSX1_114 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_29_), .Q(memory_12__1_) );
DFFPOSX1 DFFPOSX1_115 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_30_), .Q(memory_12__2_) );
DFFPOSX1 DFFPOSX1_116 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_31_), .Q(memory_12__3_) );
DFFPOSX1 DFFPOSX1_117 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_32_), .Q(memory_12__4_) );
DFFPOSX1 DFFPOSX1_118 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_33_), .Q(memory_12__5_) );
DFFPOSX1 DFFPOSX1_119 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_34_), .Q(memory_12__6_) );
DFFPOSX1 DFFPOSX1_120 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_35_), .Q(memory_12__7_) );
DFFPOSX1 DFFPOSX1_121 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_20_), .Q(memory_11__0_) );
DFFPOSX1 DFFPOSX1_122 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_21_), .Q(memory_11__1_) );
DFFPOSX1 DFFPOSX1_123 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_22_), .Q(memory_11__2_) );
DFFPOSX1 DFFPOSX1_124 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_23_), .Q(memory_11__3_) );
DFFPOSX1 DFFPOSX1_125 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_24_), .Q(memory_11__4_) );
DFFPOSX1 DFFPOSX1_126 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_25_), .Q(memory_11__5_) );
DFFPOSX1 DFFPOSX1_127 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_26_), .Q(memory_11__6_) );
DFFPOSX1 DFFPOSX1_128 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_27_), .Q(memory_11__7_) );
DFFSR DFFSR_1 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_2__0_), .Q(rd_ptr_0_), .R(_132__bF_buf3), .S(vdd) );
DFFSR DFFSR_2 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_2__1_), .Q(rd_ptr_1_), .R(_132__bF_buf2), .S(vdd) );
DFFSR DFFSR_3 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_2__2_), .Q(rd_ptr_2_), .R(_132__bF_buf1), .S(vdd) );
DFFSR DFFSR_4 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_2__3_), .Q(rd_ptr_3_), .R(_132__bF_buf0), .S(vdd) );
DFFSR DFFSR_5 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_3__0_), .Q(wr_ptr_0_), .R(_132__bF_buf3), .S(vdd) );
DFFSR DFFSR_6 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_3__1_), .Q(wr_ptr_1_), .R(_132__bF_buf2), .S(vdd) );
DFFSR DFFSR_7 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_3__2_), .Q(wr_ptr_2_), .R(_132__bF_buf1), .S(vdd) );
DFFSR DFFSR_8 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_3__3_), .Q(wr_ptr_3_), .R(_132__bF_buf0), .S(vdd) );
DFFSR DFFSR_9 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_0__0_), .Q(_568__0_), .R(_132__bF_buf3), .S(vdd) );
DFFSR DFFSR_10 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_0__1_), .Q(_568__1_), .R(_132__bF_buf2), .S(vdd) );
DFFSR DFFSR_11 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_0__2_), .Q(_568__2_), .R(_132__bF_buf1), .S(vdd) );
DFFSR DFFSR_12 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_0__3_), .Q(_568__3_), .R(_132__bF_buf0), .S(vdd) );
DFFSR DFFSR_13 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_0__4_), .Q(_568__4_), .R(_132__bF_buf3), .S(vdd) );
DFFSR DFFSR_14 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_0__5_), .Q(_568__5_), .R(_132__bF_buf2), .S(vdd) );
DFFSR DFFSR_15 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_0__6_), .Q(_568__6_), .R(_132__bF_buf1), .S(vdd) );
DFFSR DFFSR_16 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_0__7_), .Q(_568__7_), .R(_132__bF_buf0), .S(vdd) );
DFFSR DFFSR_17 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_1__0_), .Q(_570__0_), .R(_132__bF_buf3), .S(vdd) );
DFFSR DFFSR_18 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_1__1_), .Q(_570__1_), .R(_132__bF_buf2), .S(vdd) );
DFFSR DFFSR_19 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_1__2_), .Q(_570__2_), .R(_132__bF_buf1), .S(vdd) );
DFFSR DFFSR_20 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_1__3_), .Q(_570__3_), .R(_132__bF_buf0), .S(vdd) );
DFFSR DFFSR_21 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_1__4_), .Q(_570__4_), .R(_132__bF_buf3), .S(vdd) );
NOR2X1 NOR2X1_26 ( .gnd(gnd), .vdd(vdd), .A(_570__1_), .B(_570__0_), .Y(_133_) );
NOR2X1 NOR2X1_27 ( .gnd(gnd), .vdd(vdd), .A(_570__3_), .B(_570__2_), .Y(_134_) );
NAND3X1 NAND3X1_5 ( .gnd(gnd), .vdd(vdd), .A(_570__4_), .B(_133_), .C(_134_), .Y(_135_) );
INVX1 INVX1_1 ( .gnd(gnd), .vdd(vdd), .A(_135_), .Y(_571_) );
INVX2 INVX2_1 ( .gnd(gnd), .vdd(vdd), .A(_570__4_), .Y(_136_) );
NAND3X1 NAND3X1_6 ( .gnd(gnd), .vdd(vdd), .A(_136_), .B(_133_), .C(_134_), .Y(_137_) );
INVX1 INVX1_2 ( .gnd(gnd), .vdd(vdd), .A(_137_), .Y(_569_) );
INVX1 INVX1_3 ( .gnd(gnd), .vdd(vdd), .A(wr_ptr_3_), .Y(_138_) );
INVX2 INVX2_2 ( .gnd(gnd), .vdd(vdd), .A(wr_ptr_2_), .Y(_139_) );
NOR2X1 NOR2X1_28 ( .gnd(gnd), .vdd(vdd), .A(_138_), .B(_139_), .Y(_140_) );
AND2X2 AND2X2_1 ( .gnd(gnd), .vdd(vdd), .A(_135_), .B(wr_en), .Y(_141_) );
INVX2 INVX2_3 ( .gnd(gnd), .vdd(vdd), .A(wr_ptr_1_), .Y(_142_) );
INVX1 INVX1_4 ( .gnd(gnd), .vdd(vdd), .A(wr_ptr_0_), .Y(_143_) );
NOR2X1 NOR2X1_29 ( .gnd(gnd), .vdd(vdd), .A(_142_), .B(_143_), .Y(_144_) );
NAND3X1 NAND3X1_7 ( .gnd(gnd), .vdd(vdd), .A(_140_), .B(_144_), .C(_141__bF_buf0), .Y(_145_) );
NAND2X1 NAND2X1_51 ( .gnd(gnd), .vdd(vdd), .A(d_in[7]), .B(_141__bF_buf4), .Y(_146_) );
NAND2X1 NAND2X1_52 ( .gnd(gnd), .vdd(vdd), .A(memory_15__7_), .B(_145_), .Y(_147_) );
OAI21X1 OAI21X1_48 ( .gnd(gnd), .vdd(vdd), .A(_145_), .B(_146_), .C(_147_), .Y(_59_) );
NAND2X1 NAND2X1_53 ( .gnd(gnd), .vdd(vdd), .A(_133_), .B(_134_), .Y(_148_) );
OAI21X1 OAI21X1_49 ( .gnd(gnd), .vdd(vdd), .A(_148_), .B(_136_), .C(wr_en), .Y(_149_) );
AND2X2 AND2X2_2 ( .gnd(gnd), .vdd(vdd), .A(_137_), .B(rd_en), .Y(_150_) );
NAND2X1 NAND2X1_54 ( .gnd(gnd), .vdd(vdd), .A(_149_), .B(_150_), .Y(_151_) );
XNOR2X1 XNOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(_151_), .B(rd_ptr_0_bF_buf5_), .Y(_2__0_) );
OAI21X1 OAI21X1_50 ( .gnd(gnd), .vdd(vdd), .A(_148_), .B(_570__4_), .C(rd_en), .Y(_152_) );
NOR2X1 NOR2X1_30 ( .gnd(gnd), .vdd(vdd), .A(_152_), .B(_141__bF_buf3), .Y(_153_) );
AOI21X1 AOI21X1_22 ( .gnd(gnd), .vdd(vdd), .A(rd_ptr_0_bF_buf4_), .B(_153_), .C(rd_ptr_1_bF_buf3_), .Y(_154_) );
INVX8 INVX8_2 ( .gnd(gnd), .vdd(vdd), .A(rd_ptr_0_bF_buf3_), .Y(_155_) );
INVX8 INVX8_3 ( .gnd(gnd), .vdd(vdd), .A(rd_ptr_1_bF_buf2_), .Y(_156_) );
NOR2X1 NOR2X1_31 ( .gnd(gnd), .vdd(vdd), .A(_155__bF_buf5), .B(_156__bF_buf5), .Y(_157_) );
AOI21X1 AOI21X1_23 ( .gnd(gnd), .vdd(vdd), .A(_153_), .B(_157_), .C(_154_), .Y(_2__1_) );
INVX1 INVX1_5 ( .gnd(gnd), .vdd(vdd), .A(_157_), .Y(_158_) );
OAI21X1 OAI21X1_51 ( .gnd(gnd), .vdd(vdd), .A(_151_), .B(_158_), .C(rd_ptr_2_), .Y(_159_) );
INVX8 INVX8_4 ( .gnd(gnd), .vdd(vdd), .A(rd_ptr_2_), .Y(_160_) );
NAND3X1 NAND3X1_8 ( .gnd(gnd), .vdd(vdd), .A(_160__bF_buf7), .B(_157_), .C(_153_), .Y(_161_) );
NAND2X1 NAND2X1_55 ( .gnd(gnd), .vdd(vdd), .A(_159_), .B(_161_), .Y(_2__2_) );
NAND2X1 NAND2X1_56 ( .gnd(gnd), .vdd(vdd), .A(rd_ptr_2_), .B(_157_), .Y(_162_) );
XNOR2X1 XNOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(_162_), .B(rd_ptr_3_bF_buf3_), .Y(_163_) );
MUX2X1 MUX2X1_12 ( .gnd(gnd), .vdd(vdd), .A(_163_), .B(rd_ptr_3_bF_buf2_), .S(_150_), .Y(_164_) );
NAND2X1 NAND2X1_57 ( .gnd(gnd), .vdd(vdd), .A(rd_ptr_3_bF_buf1_), .B(_141__bF_buf2), .Y(_165_) );
OAI21X1 OAI21X1_52 ( .gnd(gnd), .vdd(vdd), .A(_164_), .B(_141__bF_buf1), .C(_165_), .Y(_2__3_) );
XNOR2X1 XNOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(_149_), .B(wr_ptr_0_), .Y(_3__0_) );
NOR2X1 NOR2X1_32 ( .gnd(gnd), .vdd(vdd), .A(wr_ptr_0_), .B(_142_), .Y(_166_) );
NOR2X1 NOR2X1_33 ( .gnd(gnd), .vdd(vdd), .A(wr_ptr_1_), .B(_143_), .Y(_167_) );
OAI21X1 OAI21X1_53 ( .gnd(gnd), .vdd(vdd), .A(_166_), .B(_167_), .C(_141__bF_buf0), .Y(_168_) );
OAI21X1 OAI21X1_54 ( .gnd(gnd), .vdd(vdd), .A(_142_), .B(_141__bF_buf4), .C(_168_), .Y(_3__1_) );
NAND2X1 NAND2X1_58 ( .gnd(gnd), .vdd(vdd), .A(_144_), .B(_141__bF_buf3), .Y(_169_) );
XNOR2X1 XNOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(_169_), .B(wr_ptr_2_), .Y(_3__2_) );
NOR2X1 NOR2X1_34 ( .gnd(gnd), .vdd(vdd), .A(wr_ptr_3_), .B(_139_), .Y(_170_) );
NAND3X1 NAND3X1_9 ( .gnd(gnd), .vdd(vdd), .A(_144_), .B(_170_), .C(_141__bF_buf2), .Y(_171_) );
OAI21X1 OAI21X1_55 ( .gnd(gnd), .vdd(vdd), .A(_169_), .B(_139_), .C(wr_ptr_3_), .Y(_172_) );
NAND2X1 NAND2X1_59 ( .gnd(gnd), .vdd(vdd), .A(_171__bF_buf3), .B(_172_), .Y(_3__3_) );
XNOR2X1 XNOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(_152_), .B(_570__0_), .Y(_173_) );
XNOR2X1 XNOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(_173_), .B(_149_), .Y(_1__0_) );
NOR2X1 NOR2X1_35 ( .gnd(gnd), .vdd(vdd), .A(_149_), .B(_152_), .Y(_174_) );
XOR2X1 XOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(_570__1_), .B(_570__0_), .Y(_175_) );
NAND3X1 NAND3X1_10 ( .gnd(gnd), .vdd(vdd), .A(wr_en), .B(_175_), .C(_135_), .Y(_176_) );
INVX1 INVX1_6 ( .gnd(gnd), .vdd(vdd), .A(_176_), .Y(_177_) );
INVX1 INVX1_7 ( .gnd(gnd), .vdd(vdd), .A(_570__1_), .Y(_178_) );
XNOR2X1 XNOR2X1_7 ( .gnd(gnd), .vdd(vdd), .A(_570__1_), .B(_570__0_), .Y(_179_) );
NAND3X1 NAND3X1_11 ( .gnd(gnd), .vdd(vdd), .A(rd_en), .B(_179_), .C(_137_), .Y(_180_) );
OAI21X1 OAI21X1_56 ( .gnd(gnd), .vdd(vdd), .A(_150_), .B(_178_), .C(_180_), .Y(_181_) );
AOI21X1 AOI21X1_24 ( .gnd(gnd), .vdd(vdd), .A(_149_), .B(_181_), .C(_177_), .Y(_182_) );
NAND2X1 NAND2X1_60 ( .gnd(gnd), .vdd(vdd), .A(_570__1_), .B(_174_), .Y(_183_) );
OAI21X1 OAI21X1_57 ( .gnd(gnd), .vdd(vdd), .A(_182_), .B(_174_), .C(_183_), .Y(_1__1_) );
AND2X2 AND2X2_3 ( .gnd(gnd), .vdd(vdd), .A(_570__1_), .B(_570__0_), .Y(_184_) );
NAND3X1 NAND3X1_12 ( .gnd(gnd), .vdd(vdd), .A(_184_), .B(_152_), .C(_141__bF_buf1), .Y(_185_) );
AOI21X1 AOI21X1_25 ( .gnd(gnd), .vdd(vdd), .A(_133_), .B(_153_), .C(_570__2_), .Y(_186_) );
NAND2X1 NAND2X1_61 ( .gnd(gnd), .vdd(vdd), .A(_570__2_), .B(_133_), .Y(_187_) );
OAI21X1 OAI21X1_58 ( .gnd(gnd), .vdd(vdd), .A(_152_), .B(_187_), .C(_149_), .Y(_188_) );
NAND2X1 NAND2X1_62 ( .gnd(gnd), .vdd(vdd), .A(_570__2_), .B(_184_), .Y(_189_) );
OAI21X1 OAI21X1_59 ( .gnd(gnd), .vdd(vdd), .A(_150_), .B(_189_), .C(_141__bF_buf0), .Y(_190_) );
AOI22X1 AOI22X1_1 ( .gnd(gnd), .vdd(vdd), .A(_188_), .B(_190_), .C(_186_), .D(_185_), .Y(_1__2_) );
AOI21X1 AOI21X1_26 ( .gnd(gnd), .vdd(vdd), .A(rd_en), .B(_137_), .C(_189_), .Y(_191_) );
NAND2X1 NAND2X1_63 ( .gnd(gnd), .vdd(vdd), .A(_191_), .B(_141__bF_buf4), .Y(_192_) );
INVX1 INVX1_8 ( .gnd(gnd), .vdd(vdd), .A(rd_en), .Y(_193_) );
NOR2X1 NOR2X1_36 ( .gnd(gnd), .vdd(vdd), .A(_193_), .B(_148_), .Y(_194_) );
AOI21X1 AOI21X1_27 ( .gnd(gnd), .vdd(vdd), .A(_570__4_), .B(_194_), .C(_570__3_), .Y(_195_) );
INVX1 INVX1_9 ( .gnd(gnd), .vdd(vdd), .A(_570__2_), .Y(_196_) );
NAND2X1 NAND2X1_64 ( .gnd(gnd), .vdd(vdd), .A(_196_), .B(_133_), .Y(_197_) );
OAI21X1 OAI21X1_60 ( .gnd(gnd), .vdd(vdd), .A(_151_), .B(_197_), .C(_192_), .Y(_198_) );
AOI22X1 AOI22X1_2 ( .gnd(gnd), .vdd(vdd), .A(_192_), .B(_195_), .C(_198_), .D(_570__3_), .Y(_1__3_) );
NAND3X1 NAND3X1_13 ( .gnd(gnd), .vdd(vdd), .A(_570__3_), .B(_191_), .C(_141__bF_buf3), .Y(_199_) );
NAND2X1 NAND2X1_65 ( .gnd(gnd), .vdd(vdd), .A(_194_), .B(_149_), .Y(_200_) );
NAND2X1 NAND2X1_66 ( .gnd(gnd), .vdd(vdd), .A(_570__3_), .B(_141__bF_buf2), .Y(_201_) );
OAI21X1 OAI21X1_61 ( .gnd(gnd), .vdd(vdd), .A(_201_), .B(_189_), .C(_200_), .Y(_202_) );
NOR2X1 NOR2X1_37 ( .gnd(gnd), .vdd(vdd), .A(_136_), .B(_174_), .Y(_203_) );
AOI22X1 AOI22X1_3 ( .gnd(gnd), .vdd(vdd), .A(_136_), .B(_199_), .C(_202_), .D(_203_), .Y(_1__4_) );
INVX1 INVX1_10 ( .gnd(gnd), .vdd(vdd), .A(memory_6__0_), .Y(_204_) );
OAI21X1 OAI21X1_62 ( .gnd(gnd), .vdd(vdd), .A(_160__bF_buf6), .B(_204_), .C(_155__bF_buf4), .Y(_205_) );
AOI21X1 AOI21X1_28 ( .gnd(gnd), .vdd(vdd), .A(_160__bF_buf5), .B(memory_2__0_), .C(_205_), .Y(_206_) );
INVX1 INVX1_11 ( .gnd(gnd), .vdd(vdd), .A(memory_7__0_), .Y(_207_) );
OAI21X1 OAI21X1_63 ( .gnd(gnd), .vdd(vdd), .A(_160__bF_buf4), .B(_207_), .C(rd_ptr_0_bF_buf2_), .Y(_208_) );
AOI21X1 AOI21X1_29 ( .gnd(gnd), .vdd(vdd), .A(_160__bF_buf3), .B(memory_3__0_), .C(_208_), .Y(_209_) );
OAI21X1 OAI21X1_64 ( .gnd(gnd), .vdd(vdd), .A(_206_), .B(_209_), .C(rd_ptr_1_bF_buf1_), .Y(_210_) );
INVX1 INVX1_12 ( .gnd(gnd), .vdd(vdd), .A(memory_4__0_), .Y(_211_) );
OAI21X1 OAI21X1_65 ( .gnd(gnd), .vdd(vdd), .A(_160__bF_buf2), .B(_211_), .C(_155__bF_buf3), .Y(_212_) );
AOI21X1 AOI21X1_30 ( .gnd(gnd), .vdd(vdd), .A(_160__bF_buf1), .B(memory_0__0_), .C(_212_), .Y(_213_) );
INVX1 INVX1_13 ( .gnd(gnd), .vdd(vdd), .A(memory_5__0_), .Y(_214_) );
OAI21X1 OAI21X1_66 ( .gnd(gnd), .vdd(vdd), .A(_160__bF_buf0), .B(_214_), .C(rd_ptr_0_bF_buf1_), .Y(_215_) );
AOI21X1 AOI21X1_31 ( .gnd(gnd), .vdd(vdd), .A(_160__bF_buf7), .B(memory_1__0_), .C(_215_), .Y(_216_) );
OAI21X1 OAI21X1_67 ( .gnd(gnd), .vdd(vdd), .A(_213_), .B(_216_), .C(_156__bF_buf4), .Y(_217_) );
AOI21X1 AOI21X1_32 ( .gnd(gnd), .vdd(vdd), .A(_210_), .B(_217_), .C(rd_ptr_3_bF_buf0_), .Y(_218_) );
INVX1 INVX1_14 ( .gnd(gnd), .vdd(vdd), .A(memory_14__0_), .Y(_219_) );
AOI21X1 AOI21X1_33 ( .gnd(gnd), .vdd(vdd), .A(memory_12__0_), .B(_156__bF_buf3), .C(rd_ptr_0_bF_buf0_), .Y(_220_) );
OAI21X1 OAI21X1_68 ( .gnd(gnd), .vdd(vdd), .A(_156__bF_buf2), .B(_219_), .C(_220_), .Y(_221_) );
INVX1 INVX1_15 ( .gnd(gnd), .vdd(vdd), .A(memory_15__0_), .Y(_222_) );
AOI21X1 AOI21X1_34 ( .gnd(gnd), .vdd(vdd), .A(memory_13__0_), .B(_156__bF_buf1), .C(_155__bF_buf2), .Y(_223_) );
OAI21X1 OAI21X1_69 ( .gnd(gnd), .vdd(vdd), .A(_156__bF_buf0), .B(_222_), .C(_223_), .Y(_224_) );
AOI21X1 AOI21X1_35 ( .gnd(gnd), .vdd(vdd), .A(_221_), .B(_224_), .C(_160__bF_buf6), .Y(_225_) );
INVX1 INVX1_16 ( .gnd(gnd), .vdd(vdd), .A(memory_10__0_), .Y(_226_) );
AOI21X1 AOI21X1_36 ( .gnd(gnd), .vdd(vdd), .A(memory_8__0_), .B(_156__bF_buf5), .C(rd_ptr_0_bF_buf5_), .Y(_227_) );
OAI21X1 OAI21X1_70 ( .gnd(gnd), .vdd(vdd), .A(_156__bF_buf4), .B(_226_), .C(_227_), .Y(_228_) );
INVX1 INVX1_17 ( .gnd(gnd), .vdd(vdd), .A(memory_11__0_), .Y(_229_) );
AOI21X1 AOI21X1_37 ( .gnd(gnd), .vdd(vdd), .A(memory_9__0_), .B(_156__bF_buf3), .C(_155__bF_buf1), .Y(_230_) );
OAI21X1 OAI21X1_71 ( .gnd(gnd), .vdd(vdd), .A(_156__bF_buf2), .B(_229_), .C(_230_), .Y(_231_) );
AOI21X1 AOI21X1_38 ( .gnd(gnd), .vdd(vdd), .A(_228_), .B(_231_), .C(rd_ptr_2_), .Y(_232_) );
OR2X2 OR2X2_1 ( .gnd(gnd), .vdd(vdd), .A(_225_), .B(_232_), .Y(_233_) );
AOI21X1 AOI21X1_39 ( .gnd(gnd), .vdd(vdd), .A(rd_ptr_3_bF_buf3_), .B(_233_), .C(_218_), .Y(_0__0_) );
INVX1 INVX1_18 ( .gnd(gnd), .vdd(vdd), .A(memory_6__1_), .Y(_234_) );
OAI21X1 OAI21X1_72 ( .gnd(gnd), .vdd(vdd), .A(_160__bF_buf5), .B(_234_), .C(_155__bF_buf0), .Y(_235_) );
AOI21X1 AOI21X1_40 ( .gnd(gnd), .vdd(vdd), .A(_160__bF_buf4), .B(memory_2__1_), .C(_235_), .Y(_236_) );
INVX1 INVX1_19 ( .gnd(gnd), .vdd(vdd), .A(memory_7__1_), .Y(_237_) );
OAI21X1 OAI21X1_73 ( .gnd(gnd), .vdd(vdd), .A(_160__bF_buf3), .B(_237_), .C(rd_ptr_0_bF_buf4_), .Y(_238_) );
AOI21X1 AOI21X1_41 ( .gnd(gnd), .vdd(vdd), .A(_160__bF_buf2), .B(memory_3__1_), .C(_238_), .Y(_239_) );
OAI21X1 OAI21X1_74 ( .gnd(gnd), .vdd(vdd), .A(_236_), .B(_239_), .C(rd_ptr_1_bF_buf0_), .Y(_240_) );
INVX1 INVX1_20 ( .gnd(gnd), .vdd(vdd), .A(memory_4__1_), .Y(_241_) );
OAI21X1 OAI21X1_75 ( .gnd(gnd), .vdd(vdd), .A(_160__bF_buf1), .B(_241_), .C(_155__bF_buf5), .Y(_242_) );
AOI21X1 AOI21X1_42 ( .gnd(gnd), .vdd(vdd), .A(_160__bF_buf0), .B(memory_0__1_), .C(_242_), .Y(_243_) );
INVX1 INVX1_21 ( .gnd(gnd), .vdd(vdd), .A(memory_5__1_), .Y(_244_) );
OAI21X1 OAI21X1_76 ( .gnd(gnd), .vdd(vdd), .A(_160__bF_buf7), .B(_244_), .C(rd_ptr_0_bF_buf3_), .Y(_245_) );
AOI21X1 AOI21X1_43 ( .gnd(gnd), .vdd(vdd), .A(_160__bF_buf6), .B(memory_1__1_), .C(_245_), .Y(_246_) );
OAI21X1 OAI21X1_77 ( .gnd(gnd), .vdd(vdd), .A(_243_), .B(_246_), .C(_156__bF_buf1), .Y(_247_) );
NAND2X1 NAND2X1_67 ( .gnd(gnd), .vdd(vdd), .A(_240_), .B(_247_), .Y(_248_) );
INVX1 INVX1_22 ( .gnd(gnd), .vdd(vdd), .A(memory_14__1_), .Y(_249_) );
AOI21X1 AOI21X1_44 ( .gnd(gnd), .vdd(vdd), .A(memory_12__1_), .B(_156__bF_buf0), .C(rd_ptr_0_bF_buf2_), .Y(_250_) );
OAI21X1 OAI21X1_78 ( .gnd(gnd), .vdd(vdd), .A(_156__bF_buf5), .B(_249_), .C(_250_), .Y(_251_) );
INVX1 INVX1_23 ( .gnd(gnd), .vdd(vdd), .A(memory_15__1_), .Y(_252_) );
AOI21X1 AOI21X1_45 ( .gnd(gnd), .vdd(vdd), .A(memory_13__1_), .B(_156__bF_buf4), .C(_155__bF_buf4), .Y(_253_) );
OAI21X1 OAI21X1_79 ( .gnd(gnd), .vdd(vdd), .A(_156__bF_buf3), .B(_252_), .C(_253_), .Y(_254_) );
AOI21X1 AOI21X1_46 ( .gnd(gnd), .vdd(vdd), .A(_251_), .B(_254_), .C(_160__bF_buf5), .Y(_255_) );
NOR2X1 NOR2X1_38 ( .gnd(gnd), .vdd(vdd), .A(rd_ptr_0_bF_buf1_), .B(memory_8__1_), .Y(_256_) );
OAI21X1 OAI21X1_80 ( .gnd(gnd), .vdd(vdd), .A(_155__bF_buf3), .B(memory_9__1_), .C(_156__bF_buf2), .Y(_257_) );
NOR2X1 NOR2X1_39 ( .gnd(gnd), .vdd(vdd), .A(memory_11__1_), .B(_155__bF_buf2), .Y(_258_) );
OAI21X1 OAI21X1_81 ( .gnd(gnd), .vdd(vdd), .A(rd_ptr_0_bF_buf0_), .B(memory_10__1_), .C(rd_ptr_1_bF_buf3_), .Y(_259_) );
OAI22X1 OAI22X1_1 ( .gnd(gnd), .vdd(vdd), .A(_258_), .B(_259_), .C(_257_), .D(_256_), .Y(_260_) );
OAI21X1 OAI21X1_82 ( .gnd(gnd), .vdd(vdd), .A(_260_), .B(rd_ptr_2_), .C(rd_ptr_3_bF_buf2_), .Y(_261_) );
OAI22X1 OAI22X1_2 ( .gnd(gnd), .vdd(vdd), .A(_261_), .B(_255_), .C(_248_), .D(rd_ptr_3_bF_buf1_), .Y(_0__1_) );
INVX1 INVX1_24 ( .gnd(gnd), .vdd(vdd), .A(memory_5__2_), .Y(_262_) );
AOI21X1 AOI21X1_47 ( .gnd(gnd), .vdd(vdd), .A(rd_ptr_0_bF_buf5_), .B(_262_), .C(rd_ptr_1_bF_buf2_), .Y(_263_) );
OAI21X1 OAI21X1_83 ( .gnd(gnd), .vdd(vdd), .A(rd_ptr_0_bF_buf4_), .B(memory_4__2_), .C(_263_), .Y(_264_) );
NOR2X1 NOR2X1_40 ( .gnd(gnd), .vdd(vdd), .A(memory_7__2_), .B(_155__bF_buf1), .Y(_265_) );
OAI21X1 OAI21X1_84 ( .gnd(gnd), .vdd(vdd), .A(rd_ptr_0_bF_buf3_), .B(memory_6__2_), .C(rd_ptr_1_bF_buf1_), .Y(_266_) );
OAI21X1 OAI21X1_85 ( .gnd(gnd), .vdd(vdd), .A(_265_), .B(_266_), .C(_264_), .Y(_267_) );
INVX1 INVX1_25 ( .gnd(gnd), .vdd(vdd), .A(memory_1__2_), .Y(_268_) );
AOI21X1 AOI21X1_48 ( .gnd(gnd), .vdd(vdd), .A(rd_ptr_0_bF_buf2_), .B(_268_), .C(rd_ptr_1_bF_buf0_), .Y(_269_) );
OAI21X1 OAI21X1_86 ( .gnd(gnd), .vdd(vdd), .A(rd_ptr_0_bF_buf1_), .B(memory_0__2_), .C(_269_), .Y(_270_) );
NOR2X1 NOR2X1_41 ( .gnd(gnd), .vdd(vdd), .A(memory_3__2_), .B(_155__bF_buf0), .Y(_271_) );
OAI21X1 OAI21X1_87 ( .gnd(gnd), .vdd(vdd), .A(rd_ptr_0_bF_buf0_), .B(memory_2__2_), .C(rd_ptr_1_bF_buf3_), .Y(_272_) );
OAI21X1 OAI21X1_88 ( .gnd(gnd), .vdd(vdd), .A(_271_), .B(_272_), .C(_270_), .Y(_273_) );
MUX2X1 MUX2X1_13 ( .gnd(gnd), .vdd(vdd), .A(_273_), .B(_267_), .S(_160__bF_buf4), .Y(_274_) );
NOR2X1 NOR2X1_42 ( .gnd(gnd), .vdd(vdd), .A(rd_ptr_0_bF_buf5_), .B(memory_8__2_), .Y(_275_) );
OAI21X1 OAI21X1_89 ( .gnd(gnd), .vdd(vdd), .A(_155__bF_buf5), .B(memory_9__2_), .C(_156__bF_buf1), .Y(_276_) );
NOR2X1 NOR2X1_43 ( .gnd(gnd), .vdd(vdd), .A(memory_11__2_), .B(_155__bF_buf4), .Y(_277_) );
OAI21X1 OAI21X1_90 ( .gnd(gnd), .vdd(vdd), .A(rd_ptr_0_bF_buf4_), .B(memory_10__2_), .C(rd_ptr_1_bF_buf2_), .Y(_278_) );
OAI22X1 OAI22X1_3 ( .gnd(gnd), .vdd(vdd), .A(_277_), .B(_278_), .C(_276_), .D(_275_), .Y(_279_) );
NOR2X1 NOR2X1_44 ( .gnd(gnd), .vdd(vdd), .A(rd_ptr_2_), .B(_279_), .Y(_280_) );
INVX1 INVX1_26 ( .gnd(gnd), .vdd(vdd), .A(memory_13__2_), .Y(_281_) );
AOI21X1 AOI21X1_49 ( .gnd(gnd), .vdd(vdd), .A(rd_ptr_0_bF_buf3_), .B(_281_), .C(rd_ptr_1_bF_buf1_), .Y(_282_) );
OAI21X1 OAI21X1_91 ( .gnd(gnd), .vdd(vdd), .A(rd_ptr_0_bF_buf2_), .B(memory_12__2_), .C(_282_), .Y(_283_) );
NOR2X1 NOR2X1_45 ( .gnd(gnd), .vdd(vdd), .A(memory_15__2_), .B(_155__bF_buf3), .Y(_284_) );
OAI21X1 OAI21X1_92 ( .gnd(gnd), .vdd(vdd), .A(rd_ptr_0_bF_buf1_), .B(memory_14__2_), .C(rd_ptr_1_bF_buf0_), .Y(_285_) );
OAI21X1 OAI21X1_93 ( .gnd(gnd), .vdd(vdd), .A(_284_), .B(_285_), .C(_283_), .Y(_286_) );
OAI21X1 OAI21X1_94 ( .gnd(gnd), .vdd(vdd), .A(_286_), .B(_160__bF_buf3), .C(rd_ptr_3_bF_buf0_), .Y(_287_) );
OAI22X1 OAI22X1_4 ( .gnd(gnd), .vdd(vdd), .A(_287_), .B(_280_), .C(_274_), .D(rd_ptr_3_bF_buf3_), .Y(_0__2_) );
INVX1 INVX1_27 ( .gnd(gnd), .vdd(vdd), .A(memory_6__3_), .Y(_288_) );
OAI21X1 OAI21X1_95 ( .gnd(gnd), .vdd(vdd), .A(_160__bF_buf2), .B(_288_), .C(_155__bF_buf2), .Y(_289_) );
AOI21X1 AOI21X1_50 ( .gnd(gnd), .vdd(vdd), .A(_160__bF_buf1), .B(memory_2__3_), .C(_289_), .Y(_290_) );
INVX1 INVX1_28 ( .gnd(gnd), .vdd(vdd), .A(memory_7__3_), .Y(_291_) );
OAI21X1 OAI21X1_96 ( .gnd(gnd), .vdd(vdd), .A(_160__bF_buf0), .B(_291_), .C(rd_ptr_0_bF_buf0_), .Y(_292_) );
AOI21X1 AOI21X1_51 ( .gnd(gnd), .vdd(vdd), .A(_160__bF_buf7), .B(memory_3__3_), .C(_292_), .Y(_293_) );
OAI21X1 OAI21X1_97 ( .gnd(gnd), .vdd(vdd), .A(_290_), .B(_293_), .C(rd_ptr_1_bF_buf3_), .Y(_294_) );
INVX1 INVX1_29 ( .gnd(gnd), .vdd(vdd), .A(memory_4__3_), .Y(_295_) );
OAI21X1 OAI21X1_98 ( .gnd(gnd), .vdd(vdd), .A(_160__bF_buf6), .B(_295_), .C(_155__bF_buf1), .Y(_296_) );
AOI21X1 AOI21X1_52 ( .gnd(gnd), .vdd(vdd), .A(_160__bF_buf5), .B(memory_0__3_), .C(_296_), .Y(_297_) );
INVX1 INVX1_30 ( .gnd(gnd), .vdd(vdd), .A(memory_5__3_), .Y(_298_) );
OAI21X1 OAI21X1_99 ( .gnd(gnd), .vdd(vdd), .A(_160__bF_buf4), .B(_298_), .C(rd_ptr_0_bF_buf5_), .Y(_299_) );
AOI21X1 AOI21X1_53 ( .gnd(gnd), .vdd(vdd), .A(_160__bF_buf3), .B(memory_1__3_), .C(_299_), .Y(_300_) );
OAI21X1 OAI21X1_100 ( .gnd(gnd), .vdd(vdd), .A(_297_), .B(_300_), .C(_156__bF_buf0), .Y(_301_) );
NAND2X1 NAND2X1_68 ( .gnd(gnd), .vdd(vdd), .A(_294_), .B(_301_), .Y(_302_) );
INVX1 INVX1_31 ( .gnd(gnd), .vdd(vdd), .A(memory_10__3_), .Y(_303_) );
AOI21X1 AOI21X1_54 ( .gnd(gnd), .vdd(vdd), .A(memory_8__3_), .B(_156__bF_buf5), .C(rd_ptr_0_bF_buf4_), .Y(_304_) );
OAI21X1 OAI21X1_101 ( .gnd(gnd), .vdd(vdd), .A(_156__bF_buf4), .B(_303_), .C(_304_), .Y(_305_) );
INVX1 INVX1_32 ( .gnd(gnd), .vdd(vdd), .A(memory_11__3_), .Y(_306_) );
AOI21X1 AOI21X1_55 ( .gnd(gnd), .vdd(vdd), .A(memory_9__3_), .B(_156__bF_buf3), .C(_155__bF_buf0), .Y(_307_) );
OAI21X1 OAI21X1_102 ( .gnd(gnd), .vdd(vdd), .A(_156__bF_buf2), .B(_306_), .C(_307_), .Y(_308_) );
AOI21X1 AOI21X1_56 ( .gnd(gnd), .vdd(vdd), .A(_305_), .B(_308_), .C(rd_ptr_2_), .Y(_309_) );
NOR2X1 NOR2X1_46 ( .gnd(gnd), .vdd(vdd), .A(rd_ptr_0_bF_buf3_), .B(memory_12__3_), .Y(_310_) );
OAI21X1 OAI21X1_103 ( .gnd(gnd), .vdd(vdd), .A(_155__bF_buf5), .B(memory_13__3_), .C(_156__bF_buf1), .Y(_311_) );
NOR2X1 NOR2X1_47 ( .gnd(gnd), .vdd(vdd), .A(memory_15__3_), .B(_155__bF_buf4), .Y(_312_) );
OAI21X1 OAI21X1_104 ( .gnd(gnd), .vdd(vdd), .A(rd_ptr_0_bF_buf2_), .B(memory_14__3_), .C(rd_ptr_1_bF_buf2_), .Y(_313_) );
OAI22X1 OAI22X1_5 ( .gnd(gnd), .vdd(vdd), .A(_312_), .B(_313_), .C(_311_), .D(_310_), .Y(_314_) );
OAI21X1 OAI21X1_105 ( .gnd(gnd), .vdd(vdd), .A(_314_), .B(_160__bF_buf2), .C(rd_ptr_3_bF_buf2_), .Y(_315_) );
OAI22X1 OAI22X1_6 ( .gnd(gnd), .vdd(vdd), .A(_315_), .B(_309_), .C(_302_), .D(rd_ptr_3_bF_buf1_), .Y(_0__3_) );
INVX1 INVX1_33 ( .gnd(gnd), .vdd(vdd), .A(memory_6__4_), .Y(_316_) );
OAI21X1 OAI21X1_106 ( .gnd(gnd), .vdd(vdd), .A(_160__bF_buf1), .B(_316_), .C(_155__bF_buf3), .Y(_317_) );
AOI21X1 AOI21X1_57 ( .gnd(gnd), .vdd(vdd), .A(_160__bF_buf0), .B(memory_2__4_), .C(_317_), .Y(_318_) );
INVX1 INVX1_34 ( .gnd(gnd), .vdd(vdd), .A(memory_7__4_), .Y(_319_) );
OAI21X1 OAI21X1_107 ( .gnd(gnd), .vdd(vdd), .A(_160__bF_buf7), .B(_319_), .C(rd_ptr_0_bF_buf1_), .Y(_320_) );
AOI21X1 AOI21X1_58 ( .gnd(gnd), .vdd(vdd), .A(_160__bF_buf6), .B(memory_3__4_), .C(_320_), .Y(_321_) );
OAI21X1 OAI21X1_108 ( .gnd(gnd), .vdd(vdd), .A(_318_), .B(_321_), .C(rd_ptr_1_bF_buf1_), .Y(_322_) );
INVX1 INVX1_35 ( .gnd(gnd), .vdd(vdd), .A(memory_4__4_), .Y(_323_) );
OAI21X1 OAI21X1_109 ( .gnd(gnd), .vdd(vdd), .A(_160__bF_buf5), .B(_323_), .C(_155__bF_buf2), .Y(_324_) );
AOI21X1 AOI21X1_59 ( .gnd(gnd), .vdd(vdd), .A(_160__bF_buf4), .B(memory_0__4_), .C(_324_), .Y(_325_) );
INVX1 INVX1_36 ( .gnd(gnd), .vdd(vdd), .A(memory_5__4_), .Y(_326_) );
OAI21X1 OAI21X1_110 ( .gnd(gnd), .vdd(vdd), .A(_160__bF_buf3), .B(_326_), .C(rd_ptr_0_bF_buf0_), .Y(_327_) );
AOI21X1 AOI21X1_60 ( .gnd(gnd), .vdd(vdd), .A(_160__bF_buf2), .B(memory_1__4_), .C(_327_), .Y(_328_) );
OAI21X1 OAI21X1_111 ( .gnd(gnd), .vdd(vdd), .A(_325_), .B(_328_), .C(_156__bF_buf0), .Y(_329_) );
NAND2X1 NAND2X1_69 ( .gnd(gnd), .vdd(vdd), .A(_322_), .B(_329_), .Y(_330_) );
INVX1 INVX1_37 ( .gnd(gnd), .vdd(vdd), .A(memory_10__4_), .Y(_331_) );
AOI21X1 AOI21X1_61 ( .gnd(gnd), .vdd(vdd), .A(memory_8__4_), .B(_156__bF_buf5), .C(rd_ptr_0_bF_buf5_), .Y(_332_) );
OAI21X1 OAI21X1_112 ( .gnd(gnd), .vdd(vdd), .A(_156__bF_buf4), .B(_331_), .C(_332_), .Y(_333_) );
INVX1 INVX1_38 ( .gnd(gnd), .vdd(vdd), .A(memory_11__4_), .Y(_334_) );
AOI21X1 AOI21X1_62 ( .gnd(gnd), .vdd(vdd), .A(memory_9__4_), .B(_156__bF_buf3), .C(_155__bF_buf1), .Y(_335_) );
OAI21X1 OAI21X1_113 ( .gnd(gnd), .vdd(vdd), .A(_156__bF_buf2), .B(_334_), .C(_335_), .Y(_336_) );
AOI21X1 AOI21X1_63 ( .gnd(gnd), .vdd(vdd), .A(_333_), .B(_336_), .C(rd_ptr_2_), .Y(_337_) );
NOR2X1 NOR2X1_48 ( .gnd(gnd), .vdd(vdd), .A(rd_ptr_0_bF_buf4_), .B(memory_12__4_), .Y(_338_) );
OAI21X1 OAI21X1_114 ( .gnd(gnd), .vdd(vdd), .A(_155__bF_buf0), .B(memory_13__4_), .C(_156__bF_buf1), .Y(_339_) );
NOR2X1 NOR2X1_49 ( .gnd(gnd), .vdd(vdd), .A(memory_15__4_), .B(_155__bF_buf5), .Y(_340_) );
OAI21X1 OAI21X1_115 ( .gnd(gnd), .vdd(vdd), .A(rd_ptr_0_bF_buf3_), .B(memory_14__4_), .C(rd_ptr_1_bF_buf0_), .Y(_341_) );
OAI22X1 OAI22X1_7 ( .gnd(gnd), .vdd(vdd), .A(_340_), .B(_341_), .C(_339_), .D(_338_), .Y(_342_) );
OAI21X1 OAI21X1_116 ( .gnd(gnd), .vdd(vdd), .A(_342_), .B(_160__bF_buf1), .C(rd_ptr_3_bF_buf0_), .Y(_343_) );
OAI22X1 OAI22X1_8 ( .gnd(gnd), .vdd(vdd), .A(_343_), .B(_337_), .C(_330_), .D(rd_ptr_3_bF_buf3_), .Y(_0__4_) );
INVX1 INVX1_39 ( .gnd(gnd), .vdd(vdd), .A(memory_6__5_), .Y(_344_) );
OAI21X1 OAI21X1_117 ( .gnd(gnd), .vdd(vdd), .A(_160__bF_buf0), .B(_344_), .C(_155__bF_buf4), .Y(_345_) );
AOI21X1 AOI21X1_64 ( .gnd(gnd), .vdd(vdd), .A(_160__bF_buf7), .B(memory_2__5_), .C(_345_), .Y(_346_) );
INVX1 INVX1_40 ( .gnd(gnd), .vdd(vdd), .A(memory_7__5_), .Y(_347_) );
OAI21X1 OAI21X1_118 ( .gnd(gnd), .vdd(vdd), .A(_160__bF_buf6), .B(_347_), .C(rd_ptr_0_bF_buf2_), .Y(_348_) );
AOI21X1 AOI21X1_65 ( .gnd(gnd), .vdd(vdd), .A(_160__bF_buf5), .B(memory_3__5_), .C(_348_), .Y(_349_) );
OAI21X1 OAI21X1_119 ( .gnd(gnd), .vdd(vdd), .A(_346_), .B(_349_), .C(rd_ptr_1_bF_buf3_), .Y(_350_) );
INVX1 INVX1_41 ( .gnd(gnd), .vdd(vdd), .A(memory_4__5_), .Y(_351_) );
OAI21X1 OAI21X1_120 ( .gnd(gnd), .vdd(vdd), .A(_160__bF_buf4), .B(_351_), .C(_155__bF_buf3), .Y(_352_) );
AOI21X1 AOI21X1_66 ( .gnd(gnd), .vdd(vdd), .A(_160__bF_buf3), .B(memory_0__5_), .C(_352_), .Y(_353_) );
INVX1 INVX1_42 ( .gnd(gnd), .vdd(vdd), .A(memory_5__5_), .Y(_354_) );
OAI21X1 OAI21X1_121 ( .gnd(gnd), .vdd(vdd), .A(_160__bF_buf2), .B(_354_), .C(rd_ptr_0_bF_buf1_), .Y(_355_) );
AOI21X1 AOI21X1_67 ( .gnd(gnd), .vdd(vdd), .A(_160__bF_buf1), .B(memory_1__5_), .C(_355_), .Y(_356_) );
OAI21X1 OAI21X1_122 ( .gnd(gnd), .vdd(vdd), .A(_353_), .B(_356_), .C(_156__bF_buf0), .Y(_357_) );
NAND2X1 NAND2X1_70 ( .gnd(gnd), .vdd(vdd), .A(_350_), .B(_357_), .Y(_358_) );
INVX1 INVX1_43 ( .gnd(gnd), .vdd(vdd), .A(memory_14__5_), .Y(_359_) );
AOI21X1 AOI21X1_68 ( .gnd(gnd), .vdd(vdd), .A(memory_12__5_), .B(_156__bF_buf5), .C(rd_ptr_0_bF_buf0_), .Y(_360_) );
OAI21X1 OAI21X1_123 ( .gnd(gnd), .vdd(vdd), .A(_156__bF_buf4), .B(_359_), .C(_360_), .Y(_361_) );
INVX1 INVX1_44 ( .gnd(gnd), .vdd(vdd), .A(memory_15__5_), .Y(_362_) );
AOI21X1 AOI21X1_69 ( .gnd(gnd), .vdd(vdd), .A(memory_13__5_), .B(_156__bF_buf3), .C(_155__bF_buf2), .Y(_363_) );
OAI21X1 OAI21X1_124 ( .gnd(gnd), .vdd(vdd), .A(_156__bF_buf2), .B(_362_), .C(_363_), .Y(_364_) );
AOI21X1 AOI21X1_70 ( .gnd(gnd), .vdd(vdd), .A(_361_), .B(_364_), .C(_160__bF_buf0), .Y(_365_) );
NOR2X1 NOR2X1_50 ( .gnd(gnd), .vdd(vdd), .A(rd_ptr_0_bF_buf5_), .B(memory_8__5_), .Y(_366_) );
OAI21X1 OAI21X1_125 ( .gnd(gnd), .vdd(vdd), .A(_155__bF_buf1), .B(memory_9__5_), .C(_156__bF_buf1), .Y(_367_) );
NOR2X1 NOR2X1_51 ( .gnd(gnd), .vdd(vdd), .A(memory_11__5_), .B(_155__bF_buf0), .Y(_368_) );
OAI21X1 OAI21X1_126 ( .gnd(gnd), .vdd(vdd), .A(rd_ptr_0_bF_buf4_), .B(memory_10__5_), .C(rd_ptr_1_bF_buf2_), .Y(_369_) );
OAI22X1 OAI22X1_9 ( .gnd(gnd), .vdd(vdd), .A(_368_), .B(_369_), .C(_367_), .D(_366_), .Y(_370_) );
OAI21X1 OAI21X1_127 ( .gnd(gnd), .vdd(vdd), .A(_370_), .B(rd_ptr_2_), .C(rd_ptr_3_bF_buf2_), .Y(_371_) );
OAI22X1 OAI22X1_10 ( .gnd(gnd), .vdd(vdd), .A(_371_), .B(_365_), .C(_358_), .D(rd_ptr_3_bF_buf1_), .Y(_0__5_) );
INVX1 INVX1_45 ( .gnd(gnd), .vdd(vdd), .A(memory_6__6_), .Y(_372_) );
OAI21X1 OAI21X1_128 ( .gnd(gnd), .vdd(vdd), .A(_160__bF_buf7), .B(_372_), .C(_155__bF_buf5), .Y(_373_) );
AOI21X1 AOI21X1_71 ( .gnd(gnd), .vdd(vdd), .A(_160__bF_buf6), .B(memory_2__6_), .C(_373_), .Y(_374_) );
INVX1 INVX1_46 ( .gnd(gnd), .vdd(vdd), .A(memory_7__6_), .Y(_375_) );
OAI21X1 OAI21X1_129 ( .gnd(gnd), .vdd(vdd), .A(_160__bF_buf5), .B(_375_), .C(rd_ptr_0_bF_buf3_), .Y(_376_) );
AOI21X1 AOI21X1_72 ( .gnd(gnd), .vdd(vdd), .A(_160__bF_buf4), .B(memory_3__6_), .C(_376_), .Y(_377_) );
OAI21X1 OAI21X1_130 ( .gnd(gnd), .vdd(vdd), .A(_374_), .B(_377_), .C(rd_ptr_1_bF_buf1_), .Y(_378_) );
INVX1 INVX1_47 ( .gnd(gnd), .vdd(vdd), .A(memory_4__6_), .Y(_379_) );
OAI21X1 OAI21X1_131 ( .gnd(gnd), .vdd(vdd), .A(_160__bF_buf3), .B(_379_), .C(_155__bF_buf4), .Y(_380_) );
AOI21X1 AOI21X1_73 ( .gnd(gnd), .vdd(vdd), .A(_160__bF_buf2), .B(memory_0__6_), .C(_380_), .Y(_381_) );
INVX1 INVX1_48 ( .gnd(gnd), .vdd(vdd), .A(memory_5__6_), .Y(_382_) );
OAI21X1 OAI21X1_132 ( .gnd(gnd), .vdd(vdd), .A(_160__bF_buf1), .B(_382_), .C(rd_ptr_0_bF_buf2_), .Y(_383_) );
AOI21X1 AOI21X1_74 ( .gnd(gnd), .vdd(vdd), .A(_160__bF_buf0), .B(memory_1__6_), .C(_383_), .Y(_384_) );
OAI21X1 OAI21X1_133 ( .gnd(gnd), .vdd(vdd), .A(_381_), .B(_384_), .C(_156__bF_buf0), .Y(_385_) );
NAND2X1 NAND2X1_71 ( .gnd(gnd), .vdd(vdd), .A(_378_), .B(_385_), .Y(_386_) );
INVX1 INVX1_49 ( .gnd(gnd), .vdd(vdd), .A(memory_10__6_), .Y(_387_) );
AOI21X1 AOI21X1_75 ( .gnd(gnd), .vdd(vdd), .A(memory_8__6_), .B(_156__bF_buf5), .C(rd_ptr_0_bF_buf1_), .Y(_388_) );
OAI21X1 OAI21X1_134 ( .gnd(gnd), .vdd(vdd), .A(_156__bF_buf4), .B(_387_), .C(_388_), .Y(_389_) );
INVX1 INVX1_50 ( .gnd(gnd), .vdd(vdd), .A(memory_11__6_), .Y(_390_) );
AOI21X1 AOI21X1_76 ( .gnd(gnd), .vdd(vdd), .A(memory_9__6_), .B(_156__bF_buf3), .C(_155__bF_buf3), .Y(_391_) );
OAI21X1 OAI21X1_135 ( .gnd(gnd), .vdd(vdd), .A(_156__bF_buf2), .B(_390_), .C(_391_), .Y(_392_) );
AOI21X1 AOI21X1_77 ( .gnd(gnd), .vdd(vdd), .A(_389_), .B(_392_), .C(rd_ptr_2_), .Y(_393_) );
NOR2X1 NOR2X1_52 ( .gnd(gnd), .vdd(vdd), .A(rd_ptr_0_bF_buf0_), .B(memory_12__6_), .Y(_394_) );
OAI21X1 OAI21X1_136 ( .gnd(gnd), .vdd(vdd), .A(_155__bF_buf2), .B(memory_13__6_), .C(_156__bF_buf1), .Y(_395_) );
NOR2X1 NOR2X1_53 ( .gnd(gnd), .vdd(vdd), .A(memory_15__6_), .B(_155__bF_buf1), .Y(_396_) );
OAI21X1 OAI21X1_137 ( .gnd(gnd), .vdd(vdd), .A(rd_ptr_0_bF_buf5_), .B(memory_14__6_), .C(rd_ptr_1_bF_buf0_), .Y(_397_) );
OAI22X1 OAI22X1_11 ( .gnd(gnd), .vdd(vdd), .A(_396_), .B(_397_), .C(_395_), .D(_394_), .Y(_398_) );
OAI21X1 OAI21X1_138 ( .gnd(gnd), .vdd(vdd), .A(_398_), .B(_160__bF_buf7), .C(rd_ptr_3_bF_buf0_), .Y(_399_) );
OAI22X1 OAI22X1_12 ( .gnd(gnd), .vdd(vdd), .A(_399_), .B(_393_), .C(_386_), .D(rd_ptr_3_bF_buf3_), .Y(_0__6_) );
INVX1 INVX1_51 ( .gnd(gnd), .vdd(vdd), .A(memory_6__7_), .Y(_400_) );
OAI21X1 OAI21X1_139 ( .gnd(gnd), .vdd(vdd), .A(_160__bF_buf6), .B(_400_), .C(_155__bF_buf0), .Y(_401_) );
AOI21X1 AOI21X1_78 ( .gnd(gnd), .vdd(vdd), .A(_160__bF_buf5), .B(memory_2__7_), .C(_401_), .Y(_402_) );
INVX1 INVX1_52 ( .gnd(gnd), .vdd(vdd), .A(memory_7__7_), .Y(_403_) );
OAI21X1 OAI21X1_140 ( .gnd(gnd), .vdd(vdd), .A(_160__bF_buf4), .B(_403_), .C(rd_ptr_0_bF_buf4_), .Y(_404_) );
AOI21X1 AOI21X1_79 ( .gnd(gnd), .vdd(vdd), .A(_160__bF_buf3), .B(memory_3__7_), .C(_404_), .Y(_405_) );
OAI21X1 OAI21X1_141 ( .gnd(gnd), .vdd(vdd), .A(_402_), .B(_405_), .C(rd_ptr_1_bF_buf3_), .Y(_406_) );
INVX1 INVX1_53 ( .gnd(gnd), .vdd(vdd), .A(memory_4__7_), .Y(_407_) );
OAI21X1 OAI21X1_142 ( .gnd(gnd), .vdd(vdd), .A(_160__bF_buf2), .B(_407_), .C(_155__bF_buf5), .Y(_408_) );
AOI21X1 AOI21X1_80 ( .gnd(gnd), .vdd(vdd), .A(_160__bF_buf1), .B(memory_0__7_), .C(_408_), .Y(_409_) );
INVX1 INVX1_54 ( .gnd(gnd), .vdd(vdd), .A(memory_5__7_), .Y(_410_) );
OAI21X1 OAI21X1_143 ( .gnd(gnd), .vdd(vdd), .A(_160__bF_buf0), .B(_410_), .C(rd_ptr_0_bF_buf3_), .Y(_411_) );
AOI21X1 AOI21X1_81 ( .gnd(gnd), .vdd(vdd), .A(_160__bF_buf7), .B(memory_1__7_), .C(_411_), .Y(_412_) );
OAI21X1 OAI21X1_144 ( .gnd(gnd), .vdd(vdd), .A(_409_), .B(_412_), .C(_156__bF_buf0), .Y(_413_) );
NAND2X1 NAND2X1_72 ( .gnd(gnd), .vdd(vdd), .A(_406_), .B(_413_), .Y(_414_) );
INVX1 INVX1_55 ( .gnd(gnd), .vdd(vdd), .A(memory_14__7_), .Y(_415_) );
AOI21X1 AOI21X1_82 ( .gnd(gnd), .vdd(vdd), .A(memory_12__7_), .B(_156__bF_buf5), .C(rd_ptr_0_bF_buf2_), .Y(_416_) );
OAI21X1 OAI21X1_145 ( .gnd(gnd), .vdd(vdd), .A(_156__bF_buf4), .B(_415_), .C(_416_), .Y(_417_) );
INVX1 INVX1_56 ( .gnd(gnd), .vdd(vdd), .A(memory_15__7_), .Y(_418_) );
AOI21X1 AOI21X1_83 ( .gnd(gnd), .vdd(vdd), .A(memory_13__7_), .B(_156__bF_buf3), .C(_155__bF_buf4), .Y(_419_) );
OAI21X1 OAI21X1_146 ( .gnd(gnd), .vdd(vdd), .A(_418_), .B(_156__bF_buf2), .C(_419_), .Y(_420_) );
AOI21X1 AOI21X1_84 ( .gnd(gnd), .vdd(vdd), .A(_417_), .B(_420_), .C(_160__bF_buf6), .Y(_421_) );
NOR2X1 NOR2X1_54 ( .gnd(gnd), .vdd(vdd), .A(rd_ptr_0_bF_buf1_), .B(memory_8__7_), .Y(_422_) );
OAI21X1 OAI21X1_147 ( .gnd(gnd), .vdd(vdd), .A(_155__bF_buf3), .B(memory_9__7_), .C(_156__bF_buf1), .Y(_423_) );
NOR2X1 NOR2X1_55 ( .gnd(gnd), .vdd(vdd), .A(memory_11__7_), .B(_155__bF_buf2), .Y(_424_) );
OAI21X1 OAI21X1_148 ( .gnd(gnd), .vdd(vdd), .A(rd_ptr_0_bF_buf0_), .B(memory_10__7_), .C(rd_ptr_1_bF_buf2_), .Y(_425_) );
OAI22X1 OAI22X1_13 ( .gnd(gnd), .vdd(vdd), .A(_424_), .B(_425_), .C(_423_), .D(_422_), .Y(_426_) );
OAI21X1 OAI21X1_149 ( .gnd(gnd), .vdd(vdd), .A(_426_), .B(rd_ptr_2_), .C(rd_ptr_3_bF_buf2_), .Y(_427_) );
OAI22X1 OAI22X1_14 ( .gnd(gnd), .vdd(vdd), .A(_427_), .B(_421_), .C(_414_), .D(rd_ptr_3_bF_buf1_), .Y(_0__7_) );
NOR2X1 NOR2X1_56 ( .gnd(gnd), .vdd(vdd), .A(wr_ptr_3_), .B(wr_ptr_2_), .Y(_428_) );
NOR2X1 NOR2X1_57 ( .gnd(gnd), .vdd(vdd), .A(wr_ptr_1_), .B(wr_ptr_0_), .Y(_429_) );
NAND3X1 NAND3X1_14 ( .gnd(gnd), .vdd(vdd), .A(_428_), .B(_429_), .C(_141__bF_buf1), .Y(_430_) );
NAND2X1 NAND2X1_73 ( .gnd(gnd), .vdd(vdd), .A(d_in[0]), .B(_141__bF_buf0), .Y(_431_) );
NAND2X1 NAND2X1_74 ( .gnd(gnd), .vdd(vdd), .A(memory_0__0_), .B(_430_), .Y(_432_) );
OAI21X1 OAI21X1_150 ( .gnd(gnd), .vdd(vdd), .A(_430_), .B(_431_), .C(_432_), .Y(_4_) );
NAND2X1 NAND2X1_75 ( .gnd(gnd), .vdd(vdd), .A(d_in[1]), .B(_141__bF_buf4), .Y(_433_) );
NAND2X1 NAND2X1_76 ( .gnd(gnd), .vdd(vdd), .A(memory_0__1_), .B(_430_), .Y(_434_) );
OAI21X1 OAI21X1_151 ( .gnd(gnd), .vdd(vdd), .A(_430_), .B(_433_), .C(_434_), .Y(_5_) );
NAND2X1 NAND2X1_77 ( .gnd(gnd), .vdd(vdd), .A(d_in[2]), .B(_141__bF_buf3), .Y(_435_) );
NAND2X1 NAND2X1_78 ( .gnd(gnd), .vdd(vdd), .A(memory_0__2_), .B(_430_), .Y(_436_) );
OAI21X1 OAI21X1_152 ( .gnd(gnd), .vdd(vdd), .A(_430_), .B(_435_), .C(_436_), .Y(_6_) );
NAND2X1 NAND2X1_79 ( .gnd(gnd), .vdd(vdd), .A(d_in[3]), .B(_141__bF_buf2), .Y(_437_) );
NAND2X1 NAND2X1_80 ( .gnd(gnd), .vdd(vdd), .A(memory_0__3_), .B(_430_), .Y(_438_) );
OAI21X1 OAI21X1_153 ( .gnd(gnd), .vdd(vdd), .A(_430_), .B(_437_), .C(_438_), .Y(_7_) );
NAND2X1 NAND2X1_81 ( .gnd(gnd), .vdd(vdd), .A(d_in[4]), .B(_141__bF_buf1), .Y(_439_) );
NAND2X1 NAND2X1_82 ( .gnd(gnd), .vdd(vdd), .A(memory_0__4_), .B(_430_), .Y(_440_) );
OAI21X1 OAI21X1_154 ( .gnd(gnd), .vdd(vdd), .A(_430_), .B(_439_), .C(_440_), .Y(_8_) );
NAND2X1 NAND2X1_83 ( .gnd(gnd), .vdd(vdd), .A(d_in[5]), .B(_141__bF_buf0), .Y(_441_) );
NAND2X1 NAND2X1_84 ( .gnd(gnd), .vdd(vdd), .A(memory_0__5_), .B(_430_), .Y(_442_) );
OAI21X1 OAI21X1_155 ( .gnd(gnd), .vdd(vdd), .A(_430_), .B(_441_), .C(_442_), .Y(_9_) );
NAND2X1 NAND2X1_85 ( .gnd(gnd), .vdd(vdd), .A(d_in[6]), .B(_141__bF_buf4), .Y(_443_) );
NAND2X1 NAND2X1_86 ( .gnd(gnd), .vdd(vdd), .A(memory_0__6_), .B(_430_), .Y(_444_) );
OAI21X1 OAI21X1_156 ( .gnd(gnd), .vdd(vdd), .A(_430_), .B(_443_), .C(_444_), .Y(_10_) );
NAND2X1 NAND2X1_87 ( .gnd(gnd), .vdd(vdd), .A(memory_0__7_), .B(_430_), .Y(_445_) );
OAI21X1 OAI21X1_157 ( .gnd(gnd), .vdd(vdd), .A(_146_), .B(_430_), .C(_445_), .Y(_11_) );
NAND2X1 NAND2X1_88 ( .gnd(gnd), .vdd(vdd), .A(_428_), .B(_167_), .Y(_446_) );
NOR2X1 NOR2X1_58 ( .gnd(gnd), .vdd(vdd), .A(_446_), .B(_149_), .Y(_447_) );
NOR2X1 NOR2X1_59 ( .gnd(gnd), .vdd(vdd), .A(memory_1__0_), .B(_447_), .Y(_448_) );
AOI21X1 AOI21X1_85 ( .gnd(gnd), .vdd(vdd), .A(_431_), .B(_447_), .C(_448_), .Y(_60_) );
NOR2X1 NOR2X1_60 ( .gnd(gnd), .vdd(vdd), .A(memory_1__1_), .B(_447_), .Y(_449_) );
AOI21X1 AOI21X1_86 ( .gnd(gnd), .vdd(vdd), .A(_433_), .B(_447_), .C(_449_), .Y(_61_) );
MUX2X1 MUX2X1_14 ( .gnd(gnd), .vdd(vdd), .A(_435_), .B(_268_), .S(_447_), .Y(_62_) );
NOR2X1 NOR2X1_61 ( .gnd(gnd), .vdd(vdd), .A(memory_1__3_), .B(_447_), .Y(_450_) );
AOI21X1 AOI21X1_87 ( .gnd(gnd), .vdd(vdd), .A(_437_), .B(_447_), .C(_450_), .Y(_63_) );
NOR2X1 NOR2X1_62 ( .gnd(gnd), .vdd(vdd), .A(memory_1__4_), .B(_447_), .Y(_451_) );
AOI21X1 AOI21X1_88 ( .gnd(gnd), .vdd(vdd), .A(_439_), .B(_447_), .C(_451_), .Y(_64_) );
NOR2X1 NOR2X1_63 ( .gnd(gnd), .vdd(vdd), .A(memory_1__5_), .B(_447_), .Y(_452_) );
AOI21X1 AOI21X1_89 ( .gnd(gnd), .vdd(vdd), .A(_441_), .B(_447_), .C(_452_), .Y(_65_) );
NOR2X1 NOR2X1_64 ( .gnd(gnd), .vdd(vdd), .A(memory_1__6_), .B(_447_), .Y(_453_) );
AOI21X1 AOI21X1_90 ( .gnd(gnd), .vdd(vdd), .A(_443_), .B(_447_), .C(_453_), .Y(_66_) );
NOR2X1 NOR2X1_65 ( .gnd(gnd), .vdd(vdd), .A(memory_1__7_), .B(_447_), .Y(_454_) );
AOI21X1 AOI21X1_91 ( .gnd(gnd), .vdd(vdd), .A(_146_), .B(_447_), .C(_454_), .Y(_67_) );
INVX4 INVX4_1 ( .gnd(gnd), .vdd(vdd), .A(d_in[0]), .Y(_455_) );
NAND2X1 NAND2X1_89 ( .gnd(gnd), .vdd(vdd), .A(_428_), .B(_166_), .Y(_456_) );
NOR2X1 NOR2X1_66 ( .gnd(gnd), .vdd(vdd), .A(_456_), .B(_149_), .Y(_457_) );
NOR2X1 NOR2X1_67 ( .gnd(gnd), .vdd(vdd), .A(memory_2__0_), .B(_457_), .Y(_458_) );
AOI21X1 AOI21X1_92 ( .gnd(gnd), .vdd(vdd), .A(_455_), .B(_457_), .C(_458_), .Y(_68_) );
INVX4 INVX4_2 ( .gnd(gnd), .vdd(vdd), .A(d_in[1]), .Y(_459_) );
NOR2X1 NOR2X1_68 ( .gnd(gnd), .vdd(vdd), .A(memory_2__1_), .B(_457_), .Y(_460_) );
AOI21X1 AOI21X1_93 ( .gnd(gnd), .vdd(vdd), .A(_459_), .B(_457_), .C(_460_), .Y(_69_) );
INVX4 INVX4_3 ( .gnd(gnd), .vdd(vdd), .A(d_in[2]), .Y(_461_) );
NOR2X1 NOR2X1_69 ( .gnd(gnd), .vdd(vdd), .A(memory_2__2_), .B(_457_), .Y(_462_) );
AOI21X1 AOI21X1_94 ( .gnd(gnd), .vdd(vdd), .A(_461_), .B(_457_), .C(_462_), .Y(_70_) );
INVX4 INVX4_4 ( .gnd(gnd), .vdd(vdd), .A(d_in[3]), .Y(_463_) );
NOR2X1 NOR2X1_70 ( .gnd(gnd), .vdd(vdd), .A(memory_2__3_), .B(_457_), .Y(_464_) );
AOI21X1 AOI21X1_95 ( .gnd(gnd), .vdd(vdd), .A(_463_), .B(_457_), .C(_464_), .Y(_71_) );
INVX4 INVX4_5 ( .gnd(gnd), .vdd(vdd), .A(d_in[4]), .Y(_465_) );
NOR2X1 NOR2X1_71 ( .gnd(gnd), .vdd(vdd), .A(memory_2__4_), .B(_457_), .Y(_466_) );
AOI21X1 AOI21X1_96 ( .gnd(gnd), .vdd(vdd), .A(_465_), .B(_457_), .C(_466_), .Y(_72_) );
INVX4 INVX4_6 ( .gnd(gnd), .vdd(vdd), .A(d_in[5]), .Y(_467_) );
NOR2X1 NOR2X1_72 ( .gnd(gnd), .vdd(vdd), .A(memory_2__5_), .B(_457_), .Y(_468_) );
AOI21X1 AOI21X1_97 ( .gnd(gnd), .vdd(vdd), .A(_467_), .B(_457_), .C(_468_), .Y(_73_) );
INVX4 INVX4_7 ( .gnd(gnd), .vdd(vdd), .A(d_in[6]), .Y(_469_) );
NOR2X1 NOR2X1_73 ( .gnd(gnd), .vdd(vdd), .A(memory_2__6_), .B(_457_), .Y(_470_) );
AOI21X1 AOI21X1_98 ( .gnd(gnd), .vdd(vdd), .A(_469_), .B(_457_), .C(_470_), .Y(_74_) );
INVX4 INVX4_8 ( .gnd(gnd), .vdd(vdd), .A(d_in[7]), .Y(_471_) );
NOR2X1 NOR2X1_74 ( .gnd(gnd), .vdd(vdd), .A(memory_2__7_), .B(_457_), .Y(_472_) );
AOI21X1 AOI21X1_99 ( .gnd(gnd), .vdd(vdd), .A(_471_), .B(_457_), .C(_472_), .Y(_75_) );
NAND3X1 NAND3X1_15 ( .gnd(gnd), .vdd(vdd), .A(_144_), .B(_428_), .C(_141__bF_buf3), .Y(_473_) );
NAND2X1 NAND2X1_90 ( .gnd(gnd), .vdd(vdd), .A(memory_3__0_), .B(_473_), .Y(_474_) );
OAI21X1 OAI21X1_158 ( .gnd(gnd), .vdd(vdd), .A(_431_), .B(_473_), .C(_474_), .Y(_76_) );
NAND2X1 NAND2X1_91 ( .gnd(gnd), .vdd(vdd), .A(memory_3__1_), .B(_473_), .Y(_475_) );
OAI21X1 OAI21X1_159 ( .gnd(gnd), .vdd(vdd), .A(_433_), .B(_473_), .C(_475_), .Y(_77_) );
NAND2X1 NAND2X1_92 ( .gnd(gnd), .vdd(vdd), .A(memory_3__2_), .B(_473_), .Y(_476_) );
OAI21X1 OAI21X1_160 ( .gnd(gnd), .vdd(vdd), .A(_435_), .B(_473_), .C(_476_), .Y(_78_) );
NAND2X1 NAND2X1_93 ( .gnd(gnd), .vdd(vdd), .A(memory_3__3_), .B(_473_), .Y(_477_) );
OAI21X1 OAI21X1_161 ( .gnd(gnd), .vdd(vdd), .A(_437_), .B(_473_), .C(_477_), .Y(_79_) );
NAND2X1 NAND2X1_94 ( .gnd(gnd), .vdd(vdd), .A(memory_3__4_), .B(_473_), .Y(_478_) );
OAI21X1 OAI21X1_162 ( .gnd(gnd), .vdd(vdd), .A(_439_), .B(_473_), .C(_478_), .Y(_80_) );
NAND2X1 NAND2X1_95 ( .gnd(gnd), .vdd(vdd), .A(memory_3__5_), .B(_473_), .Y(_479_) );
OAI21X1 OAI21X1_163 ( .gnd(gnd), .vdd(vdd), .A(_441_), .B(_473_), .C(_479_), .Y(_81_) );
NAND2X1 NAND2X1_96 ( .gnd(gnd), .vdd(vdd), .A(memory_3__6_), .B(_473_), .Y(_480_) );
OAI21X1 OAI21X1_164 ( .gnd(gnd), .vdd(vdd), .A(_443_), .B(_473_), .C(_480_), .Y(_82_) );
NAND2X1 NAND2X1_97 ( .gnd(gnd), .vdd(vdd), .A(memory_3__7_), .B(_473_), .Y(_481_) );
OAI21X1 OAI21X1_165 ( .gnd(gnd), .vdd(vdd), .A(_146_), .B(_473_), .C(_481_), .Y(_83_) );
NAND2X1 NAND2X1_98 ( .gnd(gnd), .vdd(vdd), .A(_429_), .B(_170_), .Y(_482_) );
NOR2X1 NOR2X1_75 ( .gnd(gnd), .vdd(vdd), .A(_482_), .B(_149_), .Y(_483_) );
MUX2X1 MUX2X1_15 ( .gnd(gnd), .vdd(vdd), .A(_455_), .B(_211_), .S(_483_), .Y(_84_) );
MUX2X1 MUX2X1_16 ( .gnd(gnd), .vdd(vdd), .A(_459_), .B(_241_), .S(_483_), .Y(_85_) );
NOR2X1 NOR2X1_76 ( .gnd(gnd), .vdd(vdd), .A(memory_4__2_), .B(_483_), .Y(_484_) );
AOI21X1 AOI21X1_100 ( .gnd(gnd), .vdd(vdd), .A(_461_), .B(_483_), .C(_484_), .Y(_86_) );
MUX2X1 MUX2X1_17 ( .gnd(gnd), .vdd(vdd), .A(_463_), .B(_295_), .S(_483_), .Y(_87_) );
MUX2X1 MUX2X1_18 ( .gnd(gnd), .vdd(vdd), .A(_465_), .B(_323_), .S(_483_), .Y(_88_) );
MUX2X1 MUX2X1_19 ( .gnd(gnd), .vdd(vdd), .A(_467_), .B(_351_), .S(_483_), .Y(_89_) );
MUX2X1 MUX2X1_20 ( .gnd(gnd), .vdd(vdd), .A(_469_), .B(_379_), .S(_483_), .Y(_90_) );
MUX2X1 MUX2X1_21 ( .gnd(gnd), .vdd(vdd), .A(_471_), .B(_407_), .S(_483_), .Y(_91_) );
NAND2X1 NAND2X1_99 ( .gnd(gnd), .vdd(vdd), .A(_167_), .B(_170_), .Y(_485_) );
NOR2X1 NOR2X1_77 ( .gnd(gnd), .vdd(vdd), .A(_485_), .B(_149_), .Y(_486_) );
MUX2X1 MUX2X1_22 ( .gnd(gnd), .vdd(vdd), .A(_431_), .B(_214_), .S(_486_), .Y(_92_) );
MUX2X1 MUX2X1_23 ( .gnd(gnd), .vdd(vdd), .A(_433_), .B(_244_), .S(_486_), .Y(_93_) );
MUX2X1 MUX2X1_24 ( .gnd(gnd), .vdd(vdd), .A(_435_), .B(_262_), .S(_486_), .Y(_94_) );
MUX2X1 MUX2X1_25 ( .gnd(gnd), .vdd(vdd), .A(_437_), .B(_298_), .S(_486_), .Y(_95_) );
MUX2X1 MUX2X1_26 ( .gnd(gnd), .vdd(vdd), .A(_439_), .B(_326_), .S(_486_), .Y(_96_) );
MUX2X1 MUX2X1_27 ( .gnd(gnd), .vdd(vdd), .A(_441_), .B(_354_), .S(_486_), .Y(_97_) );
MUX2X1 MUX2X1_28 ( .gnd(gnd), .vdd(vdd), .A(_443_), .B(_382_), .S(_486_), .Y(_98_) );
MUX2X1 MUX2X1_29 ( .gnd(gnd), .vdd(vdd), .A(_146_), .B(_410_), .S(_486_), .Y(_99_) );
NAND2X1 NAND2X1_100 ( .gnd(gnd), .vdd(vdd), .A(_166_), .B(_170_), .Y(_487_) );
NOR2X1 NOR2X1_78 ( .gnd(gnd), .vdd(vdd), .A(_487_), .B(_149_), .Y(_488_) );
endmodule
