* NGSPICE file created from fifo.ext - technology: scmos

* Black-box entry subcircuit for MUX2X1 abstract view
.subckt MUX2X1 A B S gnd Y vdd
.ends

* Black-box entry subcircuit for NAND2X1 abstract view
.subckt NAND2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for DFFSR abstract view
.subckt DFFSR Q CLK R S D gnd vdd
.ends

* Black-box entry subcircuit for OAI22X1 abstract view
.subckt OAI22X1 A B C D gnd Y vdd
.ends

* Black-box entry subcircuit for FILL abstract view
.subckt FILL gnd vdd
.ends

* Black-box entry subcircuit for OAI21X1 abstract view
.subckt OAI21X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for DFFPOSX1 abstract view
.subckt DFFPOSX1 Q CLK D gnd vdd
.ends

* Black-box entry subcircuit for BUFX4 abstract view
.subckt BUFX4 A gnd Y vdd
.ends

* Black-box entry subcircuit for INVX1 abstract view
.subckt INVX1 A gnd Y vdd
.ends

* Black-box entry subcircuit for XNOR2X1 abstract view
.subckt XNOR2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for AOI22X1 abstract view
.subckt AOI22X1 A B C D gnd Y vdd
.ends

* Black-box entry subcircuit for INVX8 abstract view
.subckt INVX8 A gnd Y vdd
.ends

* Black-box entry subcircuit for CLKBUF1 abstract view
.subckt CLKBUF1 A gnd Y vdd
.ends

* Black-box entry subcircuit for AOI21X1 abstract view
.subckt AOI21X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for NAND3X1 abstract view
.subckt NAND3X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for XOR2X1 abstract view
.subckt XOR2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for INVX4 abstract view
.subckt INVX4 A gnd Y vdd
.ends

* Black-box entry subcircuit for BUFX2 abstract view
.subckt BUFX2 A gnd Y vdd
.ends

* Black-box entry subcircuit for INVX2 abstract view
.subckt INVX2 A gnd Y vdd
.ends

* Black-box entry subcircuit for NOR2X1 abstract view
.subckt NOR2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for AND2X2 abstract view
.subckt AND2X2 A B gnd Y vdd
.ends

* Black-box entry subcircuit for OR2X2 abstract view
.subckt OR2X2 A B gnd Y vdd
.ends

.subckt fifo vdd gnd clk reset d_in[0] d_in[1] d_in[2] d_in[3] d_in[4] d_in[5] d_in[6]
+ d_in[7] wr_en rd_en full empty d_out[0] d_out[1] d_out[2] d_out[3] d_out[4] d_out[5]
+ d_out[6] d_out[7] fifo_counter[0] fifo_counter[1] fifo_counter[2] fifo_counter[3]
+ fifo_counter[4]
XMUX2X1_28 OAI21X1_7/B INVX1_48/Y NOR2X1_77/Y gnd MUX2X1_28/Y vdd MUX2X1
XMUX2X1_17 INVX4_4/Y INVX1_29/Y MUX2X1_19/S gnd MUX2X1_17/Y vdd MUX2X1
XNAND2X1_10 NOR2X1_33/Y NOR2X1_2/Y gnd NOR2X1_12/A vdd NAND2X1
XDFFSR_9 BUFX2_1/A CLKBUF1_6/Y DFFSR_9/R vdd DFFSR_9/D gnd vdd DFFSR
XNAND2X1_65 NOR2X1_36/Y NOR2X1_3/B gnd OAI21X1_61/C vdd NAND2X1
XNAND2X1_54 NOR2X1_3/B AND2X2_2/Y gnd XNOR2X1_1/A vdd NAND2X1
XNAND2X1_43 INVX1_55/A NAND3X1_4/Y gnd OAI21X1_40/C vdd NAND2X1
XNAND2X1_98 NOR2X1_57/Y NOR2X1_34/Y gnd NOR2X1_75/A vdd NAND2X1
XNAND2X1_21 NAND2X1_21/A NAND3X1_2/Y gnd OAI21X1_18/C vdd NAND2X1
XNAND2X1_76 AOI21X1_42/B NAND3X1_14/Y gnd NAND2X1_76/Y vdd NAND2X1
XNAND2X1_87 AOI21X1_80/B NAND3X1_14/Y gnd NAND2X1_87/Y vdd NAND2X1
XNAND2X1_32 NAND2X1_32/A NAND3X1_3/Y gnd OAI21X1_29/C vdd NAND2X1
XOAI22X1_3 NOR2X1_43/Y OAI22X1_3/B OAI22X1_3/C OAI22X1_3/D gnd OAI22X1_3/Y vdd OAI22X1
XFILL_11_1_0 gnd vdd FILL
XOAI21X1_19 MUX2X1_24/A NAND3X1_2/Y OAI21X1_19/C gnd OAI21X1_19/Y vdd OAI21X1
XFILL_3_2_0 gnd vdd FILL
XDFFPOSX1_125 INVX1_38/A CLKBUF1_4/Y OAI21X1_13/Y gnd vdd DFFPOSX1
XDFFPOSX1_114 NAND2X1_21/A CLKBUF1_8/Y OAI21X1_18/Y gnd vdd DFFPOSX1
XDFFPOSX1_103 INVX1_48/A CLKBUF1_7/Y MUX2X1_28/Y gnd vdd DFFPOSX1
XBUFX4_41 DFFSR_1/Q gnd BUFX4_41/Y vdd BUFX4
XBUFX4_30 INVX8_4/Y gnd BUFX4_30/Y vdd BUFX4
XINVX1_6 INVX1_6/A gnd INVX1_6/Y vdd INVX1
XXNOR2X1_6 XNOR2X1_6/A NOR2X1_3/B gnd DFFSR_17/D vdd XNOR2X1
XFILL_0_0_0 gnd vdd FILL
XFILL_16_0_0 gnd vdd FILL
XFILL_8_1_0 gnd vdd FILL
XMUX2X1_18 INVX4_5/Y INVX1_35/Y MUX2X1_19/S gnd MUX2X1_18/Y vdd MUX2X1
XMUX2X1_29 OAI21X1_8/A INVX1_54/Y NOR2X1_77/Y gnd MUX2X1_29/Y vdd MUX2X1
XNAND2X1_11 NOR2X1_32/Y NOR2X1_2/Y gnd NOR2X1_21/A vdd NAND2X1
XNAND2X1_88 NOR2X1_56/Y NOR2X1_33/Y gnd NOR2X1_58/A vdd NAND2X1
XNAND2X1_55 OAI21X1_51/Y NAND3X1_8/Y gnd DFFSR_3/D vdd NAND2X1
XAOI22X1_1 AOI22X1_1/A AOI22X1_1/B AOI22X1_1/C AOI22X1_1/D gnd DFFSR_19/D vdd AOI22X1
XNAND2X1_99 NOR2X1_33/Y NOR2X1_34/Y gnd NOR2X1_77/A vdd NAND2X1
XNAND2X1_66 DFFSR_20/Q BUFX4_8/Y gnd OAI21X1_61/A vdd NAND2X1
XNAND2X1_33 AOI21X1_69/A NAND3X1_3/Y gnd NAND2X1_33/Y vdd NAND2X1
XNAND2X1_44 INVX1_15/A NAND3X1_7/Y gnd OAI21X1_41/C vdd NAND2X1
XNAND2X1_22 OAI21X1_91/B NAND3X1_2/Y gnd OAI21X1_19/C vdd NAND2X1
XNAND2X1_77 d_in[2] BUFX4_10/Y gnd MUX2X1_24/A vdd NAND2X1
XOAI22X1_4 OAI22X1_4/A OAI22X1_4/B MUX2X1_13/Y BUFX4_34/Y gnd DFFSR_11/D vdd OAI22X1
XFILL_11_1_1 gnd vdd FILL
XFILL_3_2_1 gnd vdd FILL
XDFFPOSX1_126 NOR2X1_51/A CLKBUF1_3/Y OAI21X1_14/Y gnd vdd DFFPOSX1
XDFFPOSX1_104 INVX1_54/A CLKBUF1_9/Y MUX2X1_29/Y gnd vdd DFFPOSX1
XDFFPOSX1_115 OAI21X1_91/B CLKBUF1_9/Y OAI21X1_19/Y gnd vdd DFFPOSX1
XBUFX4_42 DFFSR_1/Q gnd BUFX4_42/Y vdd BUFX4
XBUFX4_20 INVX8_2/Y gnd BUFX4_20/Y vdd BUFX4
XBUFX4_31 INVX8_4/Y gnd BUFX4_31/Y vdd BUFX4
XXNOR2X1_7 INVX1_7/A DFFSR_17/Q gnd XNOR2X1_7/Y vdd XNOR2X1
XFILL_10_1 gnd vdd FILL
XFILL_0_0_1 gnd vdd FILL
XINVX1_7 INVX1_7/A gnd INVX1_7/Y vdd INVX1
XFILL_16_0_1 gnd vdd FILL
XFILL_8_1_1 gnd vdd FILL
XNAND2X1_89 NOR2X1_56/Y NOR2X1_32/Y gnd NOR2X1_66/A vdd NAND2X1
XAOI22X1_2 AOI22X1_2/A AOI22X1_2/B AOI22X1_2/C DFFSR_20/Q gnd DFFSR_20/D vdd AOI22X1
XMUX2X1_19 INVX4_6/Y INVX1_41/Y MUX2X1_19/S gnd MUX2X1_19/Y vdd MUX2X1
XNAND2X1_45 INVX1_23/A NAND3X1_7/Y gnd NAND2X1_45/Y vdd NAND2X1
XNAND2X1_12 INVX1_17/A NAND3X1_1/Y gnd OAI21X1_9/C vdd NAND2X1
XNAND2X1_56 DFFSR_3/Q INVX1_5/A gnd XNOR2X1_2/A vdd NAND2X1
XNAND2X1_23 NOR2X1_46/B NAND3X1_2/Y gnd OAI21X1_20/C vdd NAND2X1
XNAND2X1_78 NAND2X1_78/A NAND3X1_14/Y gnd NAND2X1_78/Y vdd NAND2X1
XNAND2X1_67 OAI21X1_74/Y OAI21X1_77/Y gnd OAI22X1_2/C vdd NAND2X1
XNAND2X1_34 NAND2X1_34/A NAND3X1_3/Y gnd NAND2X1_34/Y vdd NAND2X1
XOAI22X1_5 OAI22X1_5/A OAI22X1_5/B OAI22X1_5/C OAI22X1_5/D gnd OAI22X1_5/Y vdd OAI22X1
XDFFPOSX1_116 NOR2X1_46/B CLKBUF1_4/Y OAI21X1_20/Y gnd vdd DFFPOSX1
XDFFPOSX1_105 NAND2X1_28/A CLKBUF1_1/Y OAI21X1_25/Y gnd vdd DFFPOSX1
XDFFPOSX1_127 INVX1_50/A CLKBUF1_11/Y OAI21X1_15/Y gnd vdd DFFPOSX1
XINVX8_1 reset gnd INVX8_1/Y vdd INVX8
XBUFX4_10 BUFX4_7/A gnd BUFX4_10/Y vdd BUFX4
XBUFX4_32 INVX8_4/Y gnd BUFX4_32/Y vdd BUFX4
XBUFX4_43 DFFSR_1/Q gnd BUFX4_43/Y vdd BUFX4
XBUFX4_21 INVX8_2/Y gnd BUFX4_21/Y vdd BUFX4
XINVX1_8 rd_en gnd INVX1_8/Y vdd INVX1
XAOI22X1_3 INVX2_1/Y AOI22X1_3/B AOI22X1_3/C AOI22X1_3/D gnd DFFSR_21/D vdd AOI22X1
XOAI21X1_160 MUX2X1_24/A NAND3X1_15/Y NAND2X1_92/Y gnd DFFPOSX1_3/D vdd OAI21X1
XNAND2X1_57 BUFX4_36/Y BUFX4_9/Y gnd NAND2X1_57/Y vdd NAND2X1
XNAND2X1_35 NAND2X1_35/A NAND3X1_3/Y gnd NAND2X1_35/Y vdd NAND2X1
XNAND2X1_24 NOR2X1_48/B NAND3X1_2/Y gnd NAND2X1_24/Y vdd NAND2X1
XNAND2X1_13 NOR2X1_39/A NAND3X1_1/Y gnd NAND2X1_13/Y vdd NAND2X1
XNAND2X1_46 NOR2X1_45/A NAND3X1_7/Y gnd NAND2X1_46/Y vdd NAND2X1
XNAND2X1_79 d_in[3] BUFX4_10/Y gnd OAI21X1_4/B vdd NAND2X1
XNAND2X1_68 NAND2X1_68/A NAND2X1_68/B gnd OAI22X1_6/C vdd NAND2X1
XOAI22X1_6 OAI22X1_6/A OAI22X1_6/B OAI22X1_6/C BUFX4_36/Y gnd DFFSR_12/D vdd OAI22X1
XFILL_6_2_0 gnd vdd FILL
XFILL_14_1_0 gnd vdd FILL
XDFFPOSX1_106 AOI21X1_45/A CLKBUF1_1/Y OAI21X1_26/Y gnd vdd DFFPOSX1
XDFFPOSX1_117 NOR2X1_48/B CLKBUF1_5/Y OAI21X1_21/Y gnd vdd DFFPOSX1
XDFFPOSX1_128 NOR2X1_55/A CLKBUF1_5/Y OAI21X1_16/Y gnd vdd DFFPOSX1
XFILL_3_0_0 gnd vdd FILL
XINVX8_2 INVX8_2/A gnd INVX8_2/Y vdd INVX8
XBUFX4_11 BUFX4_7/A gnd BUFX4_11/Y vdd BUFX4
XBUFX4_44 BUFX4_45/A gnd BUFX4_44/Y vdd BUFX4
XBUFX4_33 INVX8_4/Y gnd BUFX4_33/Y vdd BUFX4
XBUFX4_22 INVX8_2/Y gnd BUFX4_22/Y vdd BUFX4
XINVX1_9 INVX1_9/A gnd INVX1_9/Y vdd INVX1
XOAI21X1_161 OAI21X1_4/B NAND3X1_15/Y NAND2X1_93/Y gnd DFFPOSX1_4/D vdd OAI21X1
XOAI21X1_150 NAND3X1_14/Y OAI21X1_9/A NAND2X1_74/Y gnd OAI21X1_150/Y vdd OAI21X1
XNAND2X1_58 NOR2X1_29/Y BUFX4_11/Y gnd XNOR2X1_4/A vdd NAND2X1
XNAND2X1_47 NOR2X1_47/A NAND3X1_7/Y gnd NAND2X1_47/Y vdd NAND2X1
XNAND2X1_69 NAND2X1_69/A NAND2X1_69/B gnd OAI22X1_8/C vdd NAND2X1
XNAND2X1_25 AOI21X1_68/A NAND3X1_2/Y gnd OAI21X1_22/C vdd NAND2X1
XNAND2X1_14 NOR2X1_43/A NAND3X1_1/Y gnd NAND2X1_14/Y vdd NAND2X1
XNAND2X1_36 INVX1_14/A NAND3X1_4/Y gnd NAND2X1_36/Y vdd NAND2X1
XOAI22X1_7 OAI22X1_7/A OAI22X1_7/B OAI22X1_7/C NOR2X1_48/Y gnd OAI22X1_7/Y vdd OAI22X1
XFILL_14_1_1 gnd vdd FILL
XFILL_6_2_1 gnd vdd FILL
XDFFPOSX1_107 INVX1_26/A CLKBUF1_9/Y OAI21X1_27/Y gnd vdd DFFPOSX1
XCLKBUF1_1 clk gnd CLKBUF1_1/Y vdd CLKBUF1
XDFFPOSX1_118 AOI21X1_68/A CLKBUF1_7/Y OAI21X1_22/Y gnd vdd DFFPOSX1
XINVX8_3 INVX8_3/A gnd BUFX4_1/A vdd INVX8
XFILL_3_0_1 gnd vdd FILL
XBUFX4_12 INVX8_1/Y gnd DFFSR_9/R vdd BUFX4
XBUFX4_45 BUFX4_45/A gnd BUFX4_45/Y vdd BUFX4
XBUFX4_34 DFFSR_4/Q gnd BUFX4_34/Y vdd BUFX4
XBUFX4_23 INVX8_2/Y gnd BUFX4_23/Y vdd BUFX4
XNAND2X1_59 BUFX4_45/Y NAND2X1_59/B gnd DFFSR_8/D vdd NAND2X1
XNAND2X1_37 INVX1_22/A NAND3X1_4/Y gnd NAND2X1_37/Y vdd NAND2X1
XOAI21X1_162 MUX2X1_26/A NAND3X1_15/Y NAND2X1_94/Y gnd DFFPOSX1_5/D vdd OAI21X1
XNAND2X1_48 NOR2X1_49/A NAND3X1_7/Y gnd OAI21X1_45/C vdd NAND2X1
XOAI21X1_140 BUFX4_31/Y INVX1_52/Y BUFX4_39/Y gnd AOI21X1_79/C vdd OAI21X1
XNAND2X1_15 INVX1_32/A NAND3X1_1/Y gnd NAND2X1_15/Y vdd NAND2X1
XOAI21X1_151 NAND3X1_14/Y OAI21X1_2/B NAND2X1_76/Y gnd DFFPOSX1_58/D vdd OAI21X1
XNAND2X1_26 NOR2X1_52/B NAND3X1_2/Y gnd OAI21X1_23/C vdd NAND2X1
XOAI22X1_8 OAI22X1_8/A OAI22X1_8/B OAI22X1_8/C BUFX4_34/Y gnd DFFSR_13/D vdd OAI22X1
XAOI21X1_90 OAI21X1_7/B NOR2X1_58/Y NOR2X1_64/Y gnd AOI21X1_90/Y vdd AOI21X1
XCLKBUF1_2 clk gnd CLKBUF1_2/Y vdd CLKBUF1
XDFFPOSX1_108 NAND2X1_31/A CLKBUF1_11/Y OAI21X1_28/Y gnd vdd DFFPOSX1
XMUX2X1_1 INVX4_1/Y MUX2X1_1/B MUX2X1_5/S gnd MUX2X1_1/Y vdd MUX2X1
XDFFPOSX1_119 NOR2X1_52/B CLKBUF1_7/Y OAI21X1_23/Y gnd vdd DFFPOSX1
XBUFX4_13 INVX8_1/Y gnd DFFSR_5/R vdd BUFX4
XDFFPOSX1_90 INVX1_22/A CLKBUF1_6/Y OAI21X1_34/Y gnd vdd DFFPOSX1
XBUFX4_35 DFFSR_4/Q gnd BUFX4_35/Y vdd BUFX4
XINVX8_4 DFFSR_3/Q gnd INVX8_4/Y vdd INVX8
XBUFX4_46 BUFX4_45/A gnd BUFX4_46/Y vdd BUFX4
XBUFX4_24 INVX8_2/Y gnd BUFX4_24/Y vdd BUFX4
XFILL_12_2_0 gnd vdd FILL
XFILL_7_1 gnd vdd FILL
XNAND3X1_1 NOR2X1_29/Y NOR2X1_2/Y BUFX4_7/Y gnd NAND3X1_1/Y vdd NAND3X1
XFILL_1_1_0 gnd vdd FILL
XFILL_17_1_0 gnd vdd FILL
XOAI21X1_163 OAI21X1_6/B NAND3X1_15/Y NAND2X1_95/Y gnd DFFPOSX1_6/D vdd OAI21X1
XNAND2X1_16 INVX1_38/A NAND3X1_1/Y gnd NAND2X1_16/Y vdd NAND2X1
XNAND2X1_27 NAND2X1_27/A NAND3X1_2/Y gnd NAND2X1_27/Y vdd NAND2X1
XFILL_9_2_0 gnd vdd FILL
XOAI21X1_152 NAND3X1_14/Y MUX2X1_24/A NAND2X1_78/Y gnd DFFPOSX1_59/D vdd OAI21X1
XNAND2X1_38 NAND2X1_38/A NAND3X1_4/Y gnd OAI21X1_35/C vdd NAND2X1
XOAI21X1_141 AOI21X1_78/Y AOI21X1_79/Y BUFX4_16/Y gnd NAND2X1_72/A vdd OAI21X1
XOAI21X1_130 AOI21X1_71/Y AOI21X1_72/Y BUFX4_18/Y gnd NAND2X1_71/A vdd OAI21X1
XNAND2X1_49 INVX1_44/A NAND3X1_7/Y gnd OAI21X1_46/C vdd NAND2X1
XOAI22X1_9 OAI22X1_9/A OAI22X1_9/B OAI22X1_9/C OAI22X1_9/D gnd OAI22X1_9/Y vdd OAI22X1
XAOI21X1_91 OAI21X1_8/A NOR2X1_58/Y NOR2X1_65/Y gnd AOI21X1_91/Y vdd AOI21X1
XAOI21X1_80 BUFX4_26/Y AOI21X1_80/B AOI21X1_80/C gnd AOI21X1_80/Y vdd AOI21X1
XCLKBUF1_3 clk gnd CLKBUF1_3/Y vdd CLKBUF1
XXOR2X1_1 INVX1_7/A DFFSR_17/Q gnd XOR2X1_1/Y vdd XOR2X1
XMUX2X1_2 INVX4_2/Y INVX1_18/Y MUX2X1_5/S gnd MUX2X1_2/Y vdd MUX2X1
XDFFPOSX1_109 NAND2X1_32/A CLKBUF1_7/Y OAI21X1_29/Y gnd vdd DFFPOSX1
XFILL_6_0_0 gnd vdd FILL
XBUFX4_14 INVX8_1/Y gnd DFFSR_4/R vdd BUFX4
XBUFX4_47 BUFX4_45/A gnd BUFX4_47/Y vdd BUFX4
XBUFX4_36 DFFSR_4/Q gnd BUFX4_36/Y vdd BUFX4
XBUFX4_25 INVX8_2/Y gnd BUFX4_25/Y vdd BUFX4
XDFFPOSX1_91 NAND2X1_38/A CLKBUF1_9/Y OAI21X1_35/Y gnd vdd DFFPOSX1
XDFFPOSX1_80 NOR2X1_11/A CLKBUF1_11/Y AOI21X1_9/Y gnd vdd DFFPOSX1
XFILL_12_2_1 gnd vdd FILL
XFILL_7_2 gnd vdd FILL
XNAND3X1_2 NAND3X1_4/A NOR2X1_57/Y BUFX4_11/Y gnd NAND3X1_2/Y vdd NAND3X1
XNAND2X1_17 NOR2X1_51/A NAND3X1_1/Y gnd OAI21X1_14/C vdd NAND2X1
XOAI21X1_120 BUFX4_28/Y INVX1_41/Y BUFX4_23/Y gnd AOI21X1_66/C vdd OAI21X1
XFILL_9_2_1 gnd vdd FILL
XNAND2X1_28 NAND2X1_28/A NAND3X1_3/Y gnd NAND2X1_28/Y vdd NAND2X1
XOAI21X1_164 OAI21X1_7/B NAND3X1_15/Y NAND2X1_96/Y gnd DFFPOSX1_7/D vdd OAI21X1
XFILL_1_1_1 gnd vdd FILL
XOAI21X1_153 NAND3X1_14/Y OAI21X1_4/B NAND2X1_80/Y gnd OAI21X1_153/Y vdd OAI21X1
XOAI21X1_142 BUFX4_27/Y INVX1_53/Y BUFX4_22/Y gnd AOI21X1_80/C vdd OAI21X1
XNAND2X1_39 NAND2X1_39/A NAND3X1_4/Y gnd OAI21X1_36/C vdd NAND2X1
XOAI21X1_131 BUFX4_31/Y INVX1_47/Y BUFX4_22/Y gnd AOI21X1_73/C vdd OAI21X1
XFILL_17_1_1 gnd vdd FILL
XAOI21X1_70 AOI21X1_70/A AOI21X1_70/B BUFX4_32/Y gnd AOI21X1_70/Y vdd AOI21X1
XAOI21X1_81 BUFX4_33/Y NOR2X1_65/A AOI21X1_81/C gnd AOI21X1_81/Y vdd AOI21X1
XAOI21X1_92 INVX4_1/Y NOR2X1_66/Y NOR2X1_67/Y gnd AOI21X1_92/Y vdd AOI21X1
XCLKBUF1_4 clk gnd CLKBUF1_4/Y vdd CLKBUF1
XFILL_6_0_1 gnd vdd FILL
XMUX2X1_3 INVX4_4/Y MUX2X1_3/B MUX2X1_5/S gnd MUX2X1_3/Y vdd MUX2X1
XDFFPOSX1_70 NOR2X1_72/A CLKBUF1_2/Y AOI21X1_97/Y gnd vdd DFFPOSX1
XBUFX4_15 INVX8_1/Y gnd DFFSR_1/R vdd BUFX4
XDFFPOSX1_81 INVX1_15/A CLKBUF1_2/Y OAI21X1_41/Y gnd vdd DFFPOSX1
XBUFX4_37 DFFSR_4/Q gnd BUFX4_37/Y vdd BUFX4
XBUFX4_26 INVX8_4/Y gnd BUFX4_26/Y vdd BUFX4
XDFFPOSX1_92 NAND2X1_39/A CLKBUF1_7/Y OAI21X1_36/Y gnd vdd DFFPOSX1
XNAND3X1_3 NAND3X1_4/A NOR2X1_33/Y BUFX4_9/Y gnd NAND3X1_3/Y vdd NAND3X1
XOAI21X1_121 BUFX4_32/Y INVX1_42/Y BUFX4_42/Y gnd AOI21X1_67/C vdd OAI21X1
XOAI21X1_165 OAI21X1_8/A NAND3X1_15/Y NAND2X1_97/Y gnd DFFPOSX1_8/D vdd OAI21X1
XOAI21X1_143 BUFX4_33/Y INVX1_54/Y INVX8_2/A gnd AOI21X1_81/C vdd OAI21X1
XOAI21X1_110 BUFX4_33/Y INVX1_36/Y BUFX4_43/Y gnd AOI21X1_60/C vdd OAI21X1
XOAI21X1_132 BUFX4_29/Y INVX1_48/Y BUFX4_41/Y gnd AOI21X1_74/C vdd OAI21X1
XOAI21X1_154 NAND3X1_14/Y MUX2X1_26/A NAND2X1_82/Y gnd DFFPOSX1_61/D vdd OAI21X1
XNAND2X1_29 AOI21X1_45/A NAND3X1_3/Y gnd NAND2X1_29/Y vdd NAND2X1
XNAND2X1_18 INVX1_50/A NAND3X1_1/Y gnd OAI21X1_15/C vdd NAND2X1
XAOI21X1_82 NAND2X1_27/A BUFX4_5/Y BUFX4_41/Y gnd AOI21X1_82/Y vdd AOI21X1
XAOI21X1_60 BUFX4_26/Y NOR2X1_62/A AOI21X1_60/C gnd AOI21X1_60/Y vdd AOI21X1
XAOI21X1_93 INVX4_2/Y NOR2X1_66/Y NOR2X1_68/Y gnd AOI21X1_93/Y vdd AOI21X1
XAOI21X1_71 BUFX4_27/Y NOR2X1_73/A AOI21X1_71/C gnd AOI21X1_71/Y vdd AOI21X1
XMUX2X1_4 INVX4_5/Y MUX2X1_4/B MUX2X1_5/S gnd MUX2X1_4/Y vdd MUX2X1
XCLKBUF1_5 clk gnd CLKBUF1_5/Y vdd CLKBUF1
XDFFPOSX1_82 INVX1_23/A CLKBUF1_4/Y OAI21X1_42/Y gnd vdd DFFPOSX1
XDFFPOSX1_71 NOR2X1_73/A CLKBUF1_1/Y AOI21X1_98/Y gnd vdd DFFPOSX1
XDFFPOSX1_60 AOI21X1_52/B CLKBUF1_7/Y OAI21X1_153/Y gnd vdd DFFPOSX1
XDFFPOSX1_93 NAND2X1_40/A CLKBUF1_9/Y OAI21X1_37/Y gnd vdd DFFPOSX1
XFILL_15_2_0 gnd vdd FILL
XBUFX4_38 DFFSR_1/Q gnd BUFX4_38/Y vdd BUFX4
XBUFX4_16 DFFSR_2/Q gnd BUFX4_16/Y vdd BUFX4
XBUFX4_27 INVX8_4/Y gnd BUFX4_27/Y vdd BUFX4
XFILL_12_0_0 gnd vdd FILL
XBUFX4_1 BUFX4_1/A gnd BUFX4_1/Y vdd BUFX4
XINVX4_1 d_in[0] gnd INVX4_1/Y vdd INVX4
XFILL_4_1_0 gnd vdd FILL
XNAND3X1_4 NAND3X1_4/A NOR2X1_32/Y BUFX4_11/Y gnd NAND3X1_4/Y vdd NAND3X1
XOAI21X1_122 AOI21X1_66/Y AOI21X1_67/Y BUFX4_4/Y gnd NAND2X1_70/B vdd OAI21X1
XOAI21X1_144 AOI21X1_80/Y AOI21X1_81/Y BUFX4_3/Y gnd NAND2X1_72/B vdd OAI21X1
XOAI21X1_100 AOI21X1_52/Y AOI21X1_53/Y BUFX4_3/Y gnd NAND2X1_68/B vdd OAI21X1
XOAI21X1_111 AOI21X1_59/Y AOI21X1_60/Y BUFX4_3/Y gnd NAND2X1_69/B vdd OAI21X1
XOAI21X1_133 AOI21X1_73/Y AOI21X1_74/Y BUFX4_3/Y gnd NAND2X1_71/B vdd OAI21X1
XOAI21X1_155 NAND3X1_14/Y OAI21X1_6/B NAND2X1_84/Y gnd DFFPOSX1_62/D vdd OAI21X1
XNAND2X1_19 NOR2X1_55/A NAND3X1_1/Y gnd OAI21X1_16/C vdd NAND2X1
XAOI21X1_61 NOR2X1_8/A BUFX4_2/Y BUFX4_38/Y gnd AOI21X1_61/Y vdd AOI21X1
XOAI21X1_1 BUFX4_44/Y OAI21X1_9/A NAND2X1_1/Y gnd OAI21X1_1/Y vdd OAI21X1
XFILL_9_0_0 gnd vdd FILL
XAOI21X1_83 NAND2X1_35/A BUFX4_5/Y BUFX4_20/Y gnd AOI21X1_83/Y vdd AOI21X1
XAOI21X1_94 INVX4_3/Y NOR2X1_66/Y NOR2X1_69/Y gnd AOI21X1_94/Y vdd AOI21X1
XAOI21X1_72 BUFX4_26/Y AOI21X1_72/B AOI21X1_72/C gnd AOI21X1_72/Y vdd AOI21X1
XAOI21X1_50 BUFX4_27/Y NOR2X1_70/A AOI21X1_50/C gnd OAI21X1_97/A vdd AOI21X1
XMUX2X1_5 INVX4_6/Y INVX1_39/Y MUX2X1_5/S gnd MUX2X1_5/Y vdd MUX2X1
XCLKBUF1_6 clk gnd CLKBUF1_6/Y vdd CLKBUF1
XFILL_15_2_1 gnd vdd FILL
XBUFX4_17 DFFSR_2/Q gnd INVX8_3/A vdd BUFX4
XBUFX4_28 INVX8_4/Y gnd BUFX4_28/Y vdd BUFX4
XDFFPOSX1_94 INVX1_43/A CLKBUF1_4/Y OAI21X1_38/Y gnd vdd DFFPOSX1
XBUFX4_39 DFFSR_1/Q gnd BUFX4_39/Y vdd BUFX4
XDFFPOSX1_83 NOR2X1_45/A CLKBUF1_9/Y OAI21X1_43/Y gnd vdd DFFPOSX1
XDFFPOSX1_50 INVX1_18/A CLKBUF1_12/Y MUX2X1_2/Y gnd vdd DFFPOSX1
XDFFPOSX1_72 NOR2X1_74/A CLKBUF1_1/Y AOI21X1_99/Y gnd vdd DFFPOSX1
XDFFPOSX1_61 AOI21X1_59/B CLKBUF1_12/Y DFFPOSX1_61/D gnd vdd DFFPOSX1
XBUFX4_2 BUFX4_1/A gnd BUFX4_2/Y vdd BUFX4
XFILL_4_1_1 gnd vdd FILL
XFILL_12_0_1 gnd vdd FILL
XINVX4_2 d_in[1] gnd INVX4_2/Y vdd INVX4
XNAND3X1_5 INVX2_1/A NAND3X1_5/B NAND3X1_5/C gnd INVX1_1/A vdd NAND3X1
XOAI21X1_112 BUFX4_2/Y INVX1_37/Y AOI21X1_61/Y gnd AOI21X1_63/A vdd OAI21X1
XOAI21X1_101 BUFX4_1/Y INVX1_31/Y AOI21X1_54/Y gnd AOI21X1_56/A vdd OAI21X1
XOAI21X1_145 BUFX4_5/Y INVX1_55/Y AOI21X1_82/Y gnd AOI21X1_84/A vdd OAI21X1
XOAI21X1_123 BUFX4_5/Y INVX1_43/Y AOI21X1_68/Y gnd AOI21X1_70/A vdd OAI21X1
XOAI21X1_134 BUFX4_2/Y INVX1_49/Y AOI21X1_75/Y gnd AOI21X1_77/A vdd OAI21X1
XOAI21X1_156 NAND3X1_14/Y OAI21X1_7/B NAND2X1_86/Y gnd OAI21X1_156/Y vdd OAI21X1
XOAI21X1_2 BUFX4_45/Y OAI21X1_2/B OAI21X1_2/C gnd OAI21X1_2/Y vdd OAI21X1
XAOI21X1_62 NOR2X1_17/A BUFX4_4/Y BUFX4_21/Y gnd AOI21X1_62/Y vdd AOI21X1
XFILL_9_0_1 gnd vdd FILL
XAOI21X1_84 AOI21X1_84/A AOI21X1_84/B BUFX4_30/Y gnd OAI22X1_14/B vdd AOI21X1
XAOI21X1_95 INVX4_4/Y NOR2X1_66/Y NOR2X1_70/Y gnd AOI21X1_95/Y vdd AOI21X1
XAOI21X1_51 BUFX4_29/Y NAND2X1_93/A OAI21X1_96/Y gnd OAI21X1_97/B vdd AOI21X1
XAOI21X1_40 BUFX4_26/Y NOR2X1_68/A AOI21X1_40/C gnd AOI21X1_40/Y vdd AOI21X1
XAOI21X1_73 BUFX4_26/Y AOI21X1_73/B AOI21X1_73/C gnd AOI21X1_73/Y vdd AOI21X1
XMUX2X1_6 INVX4_7/Y INVX1_45/Y MUX2X1_5/S gnd MUX2X1_6/Y vdd MUX2X1
XCLKBUF1_7 clk gnd CLKBUF1_7/Y vdd CLKBUF1
XDFFPOSX1_95 NAND2X1_42/A CLKBUF1_6/Y OAI21X1_39/Y gnd vdd DFFPOSX1
XDFFPOSX1_84 NOR2X1_47/A CLKBUF1_4/Y OAI21X1_44/Y gnd vdd DFFPOSX1
XDFFPOSX1_40 INVX1_52/A CLKBUF1_4/Y OAI21X1_8/Y gnd vdd DFFPOSX1
XBUFX4_18 DFFSR_2/Q gnd BUFX4_18/Y vdd BUFX4
XDFFPOSX1_73 NOR2X1_4/A CLKBUF1_10/Y AOI21X1_2/Y gnd vdd DFFPOSX1
XDFFPOSX1_51 NOR2X1_1/A CLKBUF1_10/Y AOI21X1_1/Y gnd vdd DFFPOSX1
XBUFX4_29 INVX8_4/Y gnd BUFX4_29/Y vdd BUFX4
XDFFPOSX1_62 AOI21X1_66/B CLKBUF1_12/Y DFFPOSX1_62/D gnd vdd DFFPOSX1
XBUFX4_3 BUFX4_1/A gnd BUFX4_3/Y vdd BUFX4
XINVX4_3 d_in[2] gnd INVX4_3/Y vdd INVX4
XNAND3X1_6 INVX2_1/Y NAND3X1_5/B NAND3X1_5/C gnd INVX1_2/A vdd NAND3X1
XOAI21X1_113 BUFX4_4/Y INVX1_38/Y AOI21X1_62/Y gnd AOI21X1_63/B vdd OAI21X1
XOAI21X1_124 BUFX4_5/Y INVX1_44/Y AOI21X1_69/Y gnd AOI21X1_70/B vdd OAI21X1
XOAI21X1_102 BUFX4_6/Y INVX1_32/Y AOI21X1_55/Y gnd AOI21X1_56/B vdd OAI21X1
XOAI21X1_146 INVX1_56/Y BUFX4_5/Y AOI21X1_83/Y gnd AOI21X1_84/B vdd OAI21X1
XOAI21X1_135 BUFX4_1/Y INVX1_50/Y AOI21X1_76/Y gnd AOI21X1_77/B vdd OAI21X1
XOAI21X1_157 OAI21X1_8/A NAND3X1_14/Y NAND2X1_87/Y gnd OAI21X1_157/Y vdd OAI21X1
XAOI21X1_52 BUFX4_29/Y AOI21X1_52/B OAI21X1_98/Y gnd AOI21X1_52/Y vdd AOI21X1
XAOI21X1_41 BUFX4_29/Y AOI21X1_41/B AOI21X1_41/C gnd OAI21X1_74/B vdd AOI21X1
XAOI21X1_30 BUFX4_29/Y AOI21X1_30/B AOI21X1_30/C gnd AOI21X1_30/Y vdd AOI21X1
XAOI21X1_63 AOI21X1_63/A AOI21X1_63/B DFFSR_3/Q gnd OAI22X1_8/B vdd AOI21X1
XAOI21X1_96 INVX4_5/Y NOR2X1_66/Y NOR2X1_71/Y gnd AOI21X1_96/Y vdd AOI21X1
XOAI21X1_3 BUFX4_46/Y MUX2X1_24/A OAI21X1_3/C gnd OAI21X1_3/Y vdd OAI21X1
XAOI21X1_74 BUFX4_26/Y NOR2X1_64/A AOI21X1_74/C gnd AOI21X1_74/Y vdd AOI21X1
XAOI21X1_85 OAI21X1_9/A NOR2X1_58/Y NOR2X1_59/Y gnd AOI21X1_85/Y vdd AOI21X1
XCLKBUF1_8 clk gnd CLKBUF1_8/Y vdd CLKBUF1
XFILL_10_1_0 gnd vdd FILL
XFILL_2_2_0 gnd vdd FILL
XMUX2X1_7 INVX4_8/Y INVX1_51/Y MUX2X1_5/S gnd MUX2X1_7/Y vdd MUX2X1
XDFFPOSX1_96 INVX1_55/A CLKBUF1_8/Y OAI21X1_40/Y gnd vdd DFFPOSX1
XDFFPOSX1_30 NOR2X1_24/A CLKBUF1_3/Y AOI21X1_20/Y gnd vdd DFFPOSX1
XDFFPOSX1_85 NOR2X1_49/A CLKBUF1_4/Y OAI21X1_45/Y gnd vdd DFFPOSX1
XDFFPOSX1_41 NOR2X1_13/A CLKBUF1_11/Y AOI21X1_10/Y gnd vdd DFFPOSX1
XBUFX4_19 DFFSR_2/Q gnd BUFX4_19/Y vdd BUFX4
XDFFPOSX1_74 NOR2X1_5/A CLKBUF1_12/Y AOI21X1_3/Y gnd vdd DFFPOSX1
XDFFPOSX1_63 AOI21X1_73/B CLKBUF1_12/Y OAI21X1_156/Y gnd vdd DFFPOSX1
XDFFPOSX1_52 INVX1_27/A CLKBUF1_10/Y MUX2X1_3/Y gnd vdd DFFPOSX1
XFILL_15_0_0 gnd vdd FILL
XFILL_7_1_0 gnd vdd FILL
XBUFX4_4 BUFX4_1/A gnd BUFX4_4/Y vdd BUFX4
XINVX4_4 d_in[3] gnd INVX4_4/Y vdd INVX4
XNAND3X1_7 NAND3X1_4/A NOR2X1_29/Y BUFX4_7/Y gnd NAND3X1_7/Y vdd NAND3X1
XBUFX2_1 BUFX2_1/A gnd d_out[0] vdd BUFX2
XOAI21X1_125 BUFX4_21/Y NOR2X1_18/A BUFX4_4/Y gnd OAI22X1_9/C vdd OAI21X1
XOAI21X1_103 BUFX4_21/Y NAND2X1_31/A BUFX4_2/Y gnd OAI22X1_5/C vdd OAI21X1
XOAI21X1_158 OAI21X1_9/A NAND3X1_15/Y NAND2X1_90/Y gnd DFFPOSX1_1/D vdd OAI21X1
XOAI21X1_147 BUFX4_20/Y NOR2X1_20/A BUFX4_6/Y gnd OAI22X1_13/C vdd OAI21X1
XOAI21X1_114 BUFX4_20/Y NAND2X1_32/A BUFX4_6/Y gnd OAI22X1_7/C vdd OAI21X1
XOAI21X1_136 BUFX4_20/Y NAND2X1_34/A BUFX4_6/Y gnd OAI22X1_11/C vdd OAI21X1
XAOI21X1_1 INVX4_3/Y MUX2X1_5/S NOR2X1_1/Y gnd AOI21X1_1/Y vdd AOI21X1
XINVX2_1 INVX2_1/A gnd INVX2_1/Y vdd INVX2
XAOI21X1_86 OAI21X1_2/B NOR2X1_58/Y NOR2X1_60/Y gnd AOI21X1_86/Y vdd AOI21X1
XAOI21X1_97 INVX4_6/Y NOR2X1_66/Y NOR2X1_72/Y gnd AOI21X1_97/Y vdd AOI21X1
XAOI21X1_64 BUFX4_28/Y NOR2X1_72/A AOI21X1_64/C gnd AOI21X1_64/Y vdd AOI21X1
XAOI21X1_20 INVX4_6/Y MUX2X1_9/S NOR2X1_24/Y gnd AOI21X1_20/Y vdd AOI21X1
XOAI21X1_4 BUFX4_44/Y OAI21X1_4/B OAI21X1_4/C gnd OAI21X1_4/Y vdd OAI21X1
XAOI21X1_31 BUFX4_30/Y NOR2X1_59/A OAI21X1_66/Y gnd AOI21X1_31/Y vdd AOI21X1
XAOI21X1_75 NOR2X1_10/A BUFX4_2/Y BUFX4_42/Y gnd AOI21X1_75/Y vdd AOI21X1
XAOI21X1_42 BUFX4_33/Y AOI21X1_42/B AOI21X1_42/C gnd AOI21X1_42/Y vdd AOI21X1
XAOI21X1_53 BUFX4_29/Y NOR2X1_61/A OAI21X1_99/Y gnd AOI21X1_53/Y vdd AOI21X1
XFILL_3_1 gnd vdd FILL
XFILL_10_1_1 gnd vdd FILL
XCLKBUF1_9 clk gnd CLKBUF1_9/Y vdd CLKBUF1
XFILL_2_2_1 gnd vdd FILL
XMUX2X1_8 INVX4_1/Y INVX1_16/Y MUX2X1_9/S gnd MUX2X1_8/Y vdd MUX2X1
XDFFPOSX1_97 INVX1_13/A CLKBUF1_8/Y MUX2X1_22/Y gnd vdd DFFPOSX1
XDFFPOSX1_53 INVX1_33/A CLKBUF1_1/Y MUX2X1_4/Y gnd vdd DFFPOSX1
XDFFPOSX1_31 INVX1_49/A CLKBUF1_1/Y MUX2X1_11/Y gnd vdd DFFPOSX1
XDFFPOSX1_75 NOR2X1_6/A CLKBUF1_10/Y AOI21X1_4/Y gnd vdd DFFPOSX1
XDFFPOSX1_42 NOR2X1_14/A CLKBUF1_5/Y AOI21X1_11/Y gnd vdd DFFPOSX1
XDFFPOSX1_64 AOI21X1_80/B CLKBUF1_11/Y OAI21X1_157/Y gnd vdd DFFPOSX1
XDFFPOSX1_86 INVX1_44/A CLKBUF1_7/Y OAI21X1_46/Y gnd vdd DFFPOSX1
XDFFPOSX1_20 NOR2X1_61/A CLKBUF1_7/Y AOI21X1_87/Y gnd vdd DFFPOSX1
XFILL_15_0_1 gnd vdd FILL
XFILL_7_1_1 gnd vdd FILL
XBUFX4_5 BUFX4_1/A gnd BUFX4_5/Y vdd BUFX4
XINVX4_5 d_in[4] gnd INVX4_5/Y vdd INVX4
XBUFX2_2 BUFX2_2/A gnd d_out[1] vdd BUFX2
XNAND3X1_8 BUFX4_28/Y INVX1_5/A NOR2X1_30/Y gnd NAND3X1_8/Y vdd NAND3X1
XOAI21X1_126 BUFX4_39/Y NOR2X1_24/A INVX8_3/A gnd OAI22X1_9/B vdd OAI21X1
XOAI21X1_104 BUFX4_41/Y NAND2X1_39/A INVX8_3/A gnd OAI22X1_5/B vdd OAI21X1
XOAI21X1_137 BUFX4_38/Y NAND2X1_42/A BUFX4_19/Y gnd OAI22X1_11/B vdd OAI21X1
XOAI21X1_148 BUFX4_43/Y NOR2X1_25/A INVX8_3/A gnd OAI22X1_13/B vdd OAI21X1
XOAI21X1_159 OAI21X1_2/B NAND3X1_15/Y NAND2X1_91/Y gnd DFFPOSX1_2/D vdd OAI21X1
XOAI21X1_115 INVX8_2/A NAND2X1_40/A BUFX4_19/Y gnd OAI22X1_7/B vdd OAI21X1
XINVX2_2 DFFSR_7/Q gnd INVX2_2/Y vdd INVX2
XAOI21X1_2 INVX4_1/Y NOR2X1_9/B NOR2X1_4/Y gnd AOI21X1_2/Y vdd AOI21X1
XAOI21X1_65 BUFX4_32/Y NAND2X1_95/A AOI21X1_65/C gnd AOI21X1_65/Y vdd AOI21X1
XAOI21X1_43 BUFX4_32/Y NOR2X1_60/A OAI21X1_76/Y gnd OAI21X1_77/B vdd AOI21X1
XAOI21X1_10 OAI21X1_9/A NOR2X1_12/Y NOR2X1_13/Y gnd AOI21X1_10/Y vdd AOI21X1
XAOI21X1_32 OAI21X1_64/Y OAI21X1_67/Y BUFX4_37/Y gnd AOI21X1_32/Y vdd AOI21X1
XAOI21X1_54 NOR2X1_7/A BUFX4_1/Y BUFX4_39/Y gnd AOI21X1_54/Y vdd AOI21X1
XAOI21X1_21 INVX4_8/Y MUX2X1_9/S NOR2X1_25/Y gnd AOI21X1_21/Y vdd AOI21X1
XOAI21X1_5 BUFX4_46/Y MUX2X1_26/A OAI21X1_5/C gnd OAI21X1_5/Y vdd OAI21X1
XAOI21X1_98 INVX4_7/Y NOR2X1_66/Y NOR2X1_73/Y gnd AOI21X1_98/Y vdd AOI21X1
XAOI21X1_87 OAI21X1_4/B NOR2X1_58/Y NOR2X1_61/Y gnd AOI21X1_87/Y vdd AOI21X1
XAOI21X1_76 NOR2X1_19/A BUFX4_1/Y BUFX4_22/Y gnd AOI21X1_76/Y vdd AOI21X1
XMUX2X1_9 INVX4_4/Y INVX1_31/Y MUX2X1_9/S gnd MUX2X1_9/Y vdd MUX2X1
XDFFPOSX1_54 INVX1_39/A CLKBUF1_2/Y MUX2X1_5/Y gnd vdd DFFPOSX1
XDFFPOSX1_98 INVX1_21/A CLKBUF1_8/Y MUX2X1_23/Y gnd vdd DFFPOSX1
XDFFPOSX1_76 NOR2X1_7/A CLKBUF1_1/Y AOI21X1_5/Y gnd vdd DFFPOSX1
XDFFPOSX1_32 NOR2X1_25/A CLKBUF1_11/Y AOI21X1_21/Y gnd vdd DFFPOSX1
XDFFPOSX1_43 NOR2X1_15/A CLKBUF1_12/Y AOI21X1_12/Y gnd vdd DFFPOSX1
XDFFPOSX1_21 NOR2X1_62/A CLKBUF1_5/Y AOI21X1_88/Y gnd vdd DFFPOSX1
XDFFPOSX1_87 NOR2X1_53/A CLKBUF1_5/Y OAI21X1_47/Y gnd vdd DFFPOSX1
XDFFPOSX1_65 NOR2X1_67/A CLKBUF1_10/Y AOI21X1_92/Y gnd vdd DFFPOSX1
XDFFPOSX1_10 INVX1_20/A CLKBUF1_12/Y MUX2X1_16/Y gnd vdd DFFPOSX1
XINVX4_6 d_in[5] gnd INVX4_6/Y vdd INVX4
XBUFX4_6 BUFX4_1/A gnd BUFX4_6/Y vdd BUFX4
XBUFX2_3 BUFX2_3/A gnd d_out[2] vdd BUFX2
XNAND3X1_9 NOR2X1_29/Y NOR2X1_34/Y BUFX4_9/Y gnd BUFX4_45/A vdd NAND3X1
XOAI21X1_127 OAI22X1_9/Y DFFSR_3/Q BUFX4_35/Y gnd OAI22X1_10/A vdd OAI21X1
XOAI21X1_105 OAI22X1_5/Y BUFX4_31/Y BUFX4_35/Y gnd OAI22X1_6/A vdd OAI21X1
XOAI21X1_149 OAI22X1_13/Y DFFSR_3/Q BUFX4_35/Y gnd OAI22X1_14/A vdd OAI21X1
XOAI21X1_116 OAI22X1_7/Y BUFX4_30/Y BUFX4_37/Y gnd OAI22X1_8/A vdd OAI21X1
XOAI21X1_138 OAI22X1_11/Y BUFX4_30/Y BUFX4_37/Y gnd OAI22X1_12/A vdd OAI21X1
XINVX2_3 DFFSR_6/Q gnd INVX2_3/Y vdd INVX2
XNAND2X1_100 NOR2X1_32/Y NOR2X1_34/Y gnd NOR2X1_78/A vdd NAND2X1
XAOI21X1_3 INVX4_2/Y NOR2X1_9/B NOR2X1_5/Y gnd AOI21X1_3/Y vdd AOI21X1
XNOR2X1_1 NOR2X1_1/A MUX2X1_5/S gnd NOR2X1_1/Y vdd NOR2X1
XBUFX2_10 DFFSR_17/Q gnd fifo_counter[0] vdd BUFX2
XOAI21X1_6 BUFX4_44/Y OAI21X1_6/B OAI21X1_6/C gnd OAI21X1_6/Y vdd OAI21X1
XAOI21X1_66 BUFX4_28/Y AOI21X1_66/B AOI21X1_66/C gnd AOI21X1_66/Y vdd AOI21X1
XAOI21X1_44 NAND2X1_21/A BUFX4_4/Y BUFX4_41/Y gnd AOI21X1_44/Y vdd AOI21X1
XAOI21X1_22 BUFX4_39/Y NOR2X1_30/Y BUFX4_16/Y gnd AOI21X1_22/Y vdd AOI21X1
XAOI21X1_55 NOR2X1_16/A BUFX4_6/Y BUFX4_20/Y gnd AOI21X1_55/Y vdd AOI21X1
XAOI21X1_77 AOI21X1_77/A AOI21X1_77/B DFFSR_3/Q gnd OAI22X1_12/B vdd AOI21X1
XAOI21X1_11 OAI21X1_2/B NOR2X1_12/Y NOR2X1_14/Y gnd AOI21X1_11/Y vdd AOI21X1
XAOI21X1_88 MUX2X1_26/A NOR2X1_58/Y NOR2X1_62/Y gnd AOI21X1_88/Y vdd AOI21X1
XAOI21X1_33 AOI21X1_33/A BUFX4_3/Y BUFX4_43/Y gnd AOI21X1_33/Y vdd AOI21X1
XFILL_5_2_0 gnd vdd FILL
XAOI21X1_99 INVX4_8/Y NOR2X1_66/Y NOR2X1_74/Y gnd AOI21X1_99/Y vdd AOI21X1
XFILL_13_1_0 gnd vdd FILL
XDFFPOSX1_11 NOR2X1_76/A CLKBUF1_10/Y DFFPOSX1_11/D gnd vdd DFFPOSX1
XDFFPOSX1_22 NOR2X1_63/A CLKBUF1_8/Y AOI21X1_89/Y gnd vdd DFFPOSX1
XDFFPOSX1_33 INVX1_11/A CLKBUF1_8/Y OAI21X1_1/Y gnd vdd DFFPOSX1
XDFFPOSX1_77 NOR2X1_8/A CLKBUF1_3/Y AOI21X1_6/Y gnd vdd DFFPOSX1
XDFFPOSX1_55 INVX1_45/A CLKBUF1_1/Y MUX2X1_6/Y gnd vdd DFFPOSX1
XDFFPOSX1_44 NOR2X1_16/A CLKBUF1_4/Y AOI21X1_13/Y gnd vdd DFFPOSX1
XFILL_2_0_0 gnd vdd FILL
XDFFPOSX1_66 NOR2X1_68/A CLKBUF1_12/Y AOI21X1_93/Y gnd vdd DFFPOSX1
XDFFPOSX1_99 INVX1_24/A CLKBUF1_12/Y MUX2X1_24/Y gnd vdd DFFPOSX1
XDFFPOSX1_88 INVX1_56/A CLKBUF1_9/Y OAI21X1_48/Y gnd vdd DFFPOSX1
XBUFX4_7 BUFX4_7/A gnd BUFX4_7/Y vdd BUFX4
XFILL_13_1 gnd vdd FILL
XINVX4_7 d_in[6] gnd INVX4_7/Y vdd INVX4
XOAI21X1_117 BUFX4_28/Y INVX1_39/Y BUFX4_23/Y gnd AOI21X1_64/C vdd OAI21X1
XOAI21X1_106 BUFX4_28/Y MUX2X1_4/B BUFX4_23/Y gnd AOI21X1_57/C vdd OAI21X1
XOAI21X1_128 BUFX4_27/Y INVX1_45/Y BUFX4_22/Y gnd AOI21X1_71/C vdd OAI21X1
XBUFX2_4 BUFX2_4/A gnd d_out[3] vdd BUFX2
XAOI21X1_4 INVX4_3/Y NOR2X1_9/B NOR2X1_6/Y gnd AOI21X1_4/Y vdd AOI21X1
XOAI21X1_139 BUFX4_27/Y INVX1_51/Y BUFX4_22/Y gnd AOI21X1_78/C vdd OAI21X1
XNOR2X1_2 DFFSR_7/Q INVX1_3/Y gnd NOR2X1_2/Y vdd NOR2X1
XBUFX2_11 INVX1_7/A gnd fifo_counter[1] vdd BUFX2
XAOI21X1_89 OAI21X1_6/B NOR2X1_58/Y NOR2X1_63/Y gnd AOI21X1_89/Y vdd AOI21X1
XAOI21X1_67 BUFX4_32/Y NOR2X1_63/A AOI21X1_67/C gnd AOI21X1_67/Y vdd AOI21X1
XAOI21X1_23 NOR2X1_30/Y INVX1_5/A AOI21X1_22/Y gnd DFFSR_2/D vdd AOI21X1
XOAI21X1_7 BUFX4_47/Y OAI21X1_7/B NAND2X1_7/Y gnd OAI21X1_7/Y vdd OAI21X1
XAOI21X1_45 AOI21X1_45/A BUFX4_4/Y BUFX4_21/Y gnd AOI21X1_45/Y vdd AOI21X1
XAOI21X1_34 NAND2X1_28/A BUFX4_1/Y BUFX4_23/Y gnd OAI21X1_69/C vdd AOI21X1
XAOI21X1_56 AOI21X1_56/A AOI21X1_56/B DFFSR_3/Q gnd OAI22X1_6/B vdd AOI21X1
XAOI21X1_12 MUX2X1_24/A NOR2X1_12/Y NOR2X1_15/Y gnd AOI21X1_12/Y vdd AOI21X1
XAOI21X1_78 BUFX4_27/Y NOR2X1_74/A AOI21X1_78/C gnd AOI21X1_78/Y vdd AOI21X1
XFILL_13_1_1 gnd vdd FILL
XFILL_5_2_1 gnd vdd FILL
XFILL_1_1 gnd vdd FILL
XDFFPOSX1_45 NOR2X1_17/A CLKBUF1_6/Y AOI21X1_14/Y gnd vdd DFFPOSX1
XDFFPOSX1_34 INVX1_19/A CLKBUF1_3/Y OAI21X1_2/Y gnd vdd DFFPOSX1
XDFFPOSX1_78 NOR2X1_9/A CLKBUF1_3/Y AOI21X1_7/Y gnd vdd DFFPOSX1
XFILL_2_0_1 gnd vdd FILL
XDFFPOSX1_67 NOR2X1_69/A CLKBUF1_10/Y AOI21X1_94/Y gnd vdd DFFPOSX1
XDFFPOSX1_23 NOR2X1_64/A CLKBUF1_11/Y AOI21X1_90/Y gnd vdd DFFPOSX1
XDFFPOSX1_56 INVX1_51/A CLKBUF1_10/Y MUX2X1_7/Y gnd vdd DFFPOSX1
XDFFPOSX1_89 INVX1_14/A CLKBUF1_11/Y OAI21X1_33/Y gnd vdd DFFPOSX1
XDFFPOSX1_12 INVX1_29/A CLKBUF1_1/Y MUX2X1_17/Y gnd vdd DFFPOSX1
XBUFX4_8 BUFX4_7/A gnd BUFX4_8/Y vdd BUFX4
XINVX4_8 d_in[7] gnd INVX4_8/Y vdd INVX4
XBUFX2_5 BUFX2_5/A gnd d_out[4] vdd BUFX2
XOAI21X1_118 BUFX4_32/Y INVX1_40/Y BUFX4_41/Y gnd AOI21X1_65/C vdd OAI21X1
XOAI21X1_129 BUFX4_31/Y INVX1_46/Y INVX8_2/A gnd AOI21X1_72/C vdd OAI21X1
XOAI21X1_107 BUFX4_33/Y INVX1_34/Y BUFX4_42/Y gnd AOI21X1_58/C vdd OAI21X1
XAOI21X1_5 INVX4_4/Y NOR2X1_9/B NOR2X1_7/Y gnd AOI21X1_5/Y vdd AOI21X1
XBUFX2_12 INVX1_9/A gnd fifo_counter[2] vdd BUFX2
XAOI21X1_24 NOR2X1_3/B AOI21X1_24/B INVX1_6/Y gnd OAI21X1_57/A vdd AOI21X1
XNOR2X1_3 NOR2X1_3/A NOR2X1_3/B gnd NOR2X1_9/B vdd NOR2X1
XAOI21X1_46 AOI21X1_46/A AOI21X1_46/B BUFX4_32/Y gnd OAI22X1_2/B vdd AOI21X1
XAOI21X1_57 BUFX4_28/Y NOR2X1_71/A AOI21X1_57/C gnd AOI21X1_57/Y vdd AOI21X1
XAOI21X1_35 OAI21X1_68/Y AOI21X1_35/B BUFX4_31/Y gnd OR2X2_1/A vdd AOI21X1
XAOI21X1_68 AOI21X1_68/A BUFX4_5/Y BUFX4_43/Y gnd AOI21X1_68/Y vdd AOI21X1
XAOI21X1_13 OAI21X1_4/B NOR2X1_12/Y NOR2X1_16/Y gnd AOI21X1_13/Y vdd AOI21X1
XOAI22X1_10 OAI22X1_10/A AOI21X1_70/Y OAI22X1_10/C BUFX4_36/Y gnd DFFSR_14/D vdd OAI22X1
XOAI21X1_8 OAI21X1_8/A BUFX4_47/Y NAND2X1_8/Y gnd OAI21X1_8/Y vdd OAI21X1
XAOI21X1_79 BUFX4_31/Y DFFPOSX1_8/Q AOI21X1_79/C gnd AOI21X1_79/Y vdd AOI21X1
XDFFPOSX1_46 NOR2X1_18/A CLKBUF1_6/Y AOI21X1_15/Y gnd vdd DFFPOSX1
XDFFPOSX1_13 INVX1_35/A CLKBUF1_1/Y MUX2X1_18/Y gnd vdd DFFPOSX1
XDFFPOSX1_79 NOR2X1_10/A CLKBUF1_11/Y AOI21X1_8/Y gnd vdd DFFPOSX1
XDFFPOSX1_68 NOR2X1_70/A CLKBUF1_1/Y AOI21X1_95/Y gnd vdd DFFPOSX1
XDFFPOSX1_24 NOR2X1_65/A CLKBUF1_9/Y AOI21X1_91/Y gnd vdd DFFPOSX1
XDFFPOSX1_35 NOR2X1_40/A CLKBUF1_9/Y OAI21X1_3/Y gnd vdd DFFPOSX1
XDFFPOSX1_57 AOI21X1_30/B CLKBUF1_7/Y OAI21X1_150/Y gnd vdd DFFPOSX1
XAOI21X1_100 INVX4_3/Y MUX2X1_19/S NOR2X1_76/Y gnd DFFPOSX1_11/D vdd AOI21X1
XFILL_11_2_0 gnd vdd FILL
XBUFX4_9 BUFX4_7/A gnd BUFX4_9/Y vdd BUFX4
XBUFX2_6 BUFX2_6/A gnd d_out[5] vdd BUFX2
XOAI21X1_119 AOI21X1_64/Y AOI21X1_65/Y BUFX4_16/Y gnd NAND2X1_70/A vdd OAI21X1
XNAND2X1_1 INVX1_11/A BUFX4_44/Y gnd NAND2X1_1/Y vdd NAND2X1
XOAI21X1_108 AOI21X1_57/Y AOI21X1_58/Y BUFX4_18/Y gnd NAND2X1_69/A vdd OAI21X1
XFILL_16_1_0 gnd vdd FILL
XAOI21X1_6 INVX4_5/Y NOR2X1_9/B NOR2X1_8/Y gnd AOI21X1_6/Y vdd AOI21X1
XDFFPOSX1_1 AOI21X1_29/B CLKBUF1_4/Y DFFPOSX1_1/D gnd vdd DFFPOSX1
XFILL_8_2_0 gnd vdd FILL
XBUFX2_13 DFFSR_20/Q gnd fifo_counter[3] vdd BUFX2
XFILL_0_1_0 gnd vdd FILL
XNOR2X1_4 NOR2X1_4/A NOR2X1_9/B gnd NOR2X1_4/Y vdd NOR2X1
XAOI21X1_14 MUX2X1_26/A NOR2X1_12/Y NOR2X1_17/Y gnd AOI21X1_14/Y vdd AOI21X1
XAOI21X1_25 NAND3X1_5/B NOR2X1_30/Y INVX1_9/A gnd AOI22X1_1/C vdd AOI21X1
XOAI21X1_9 OAI21X1_9/A NAND3X1_1/Y OAI21X1_9/C gnd OAI21X1_9/Y vdd OAI21X1
XAOI21X1_69 AOI21X1_69/A BUFX4_5/Y BUFX4_20/Y gnd AOI21X1_69/Y vdd AOI21X1
XAOI21X1_58 BUFX4_31/Y AOI21X1_58/B AOI21X1_58/C gnd AOI21X1_58/Y vdd AOI21X1
XAOI21X1_36 NOR2X1_4/A BUFX4_1/Y BUFX4_38/Y gnd AOI21X1_36/Y vdd AOI21X1
XAOI21X1_47 BUFX4_38/Y INVX1_24/Y INVX8_3/A gnd OAI21X1_83/C vdd AOI21X1
XOAI22X1_11 NOR2X1_53/Y OAI22X1_11/B OAI22X1_11/C NOR2X1_52/Y gnd OAI22X1_11/Y vdd
+ OAI22X1
XFILL_5_0_0 gnd vdd FILL
XDFFPOSX1_14 INVX1_41/A CLKBUF1_2/Y MUX2X1_19/Y gnd vdd DFFPOSX1
XDFFPOSX1_36 INVX1_28/A CLKBUF1_4/Y OAI21X1_4/Y gnd vdd DFFPOSX1
XDFFPOSX1_69 NOR2X1_71/A CLKBUF1_3/Y AOI21X1_96/Y gnd vdd DFFPOSX1
XDFFPOSX1_25 INVX1_16/A CLKBUF1_10/Y MUX2X1_8/Y gnd vdd DFFPOSX1
XDFFPOSX1_58 AOI21X1_42/B CLKBUF1_9/Y DFFPOSX1_58/D gnd vdd DFFPOSX1
XDFFPOSX1_47 NOR2X1_19/A CLKBUF1_12/Y AOI21X1_16/Y gnd vdd DFFPOSX1
XFILL_11_2_1 gnd vdd FILL
XBUFX2_7 BUFX2_7/A gnd d_out[6] vdd BUFX2
XFILL_11_1 gnd vdd FILL
XOAI21X1_109 BUFX4_28/Y INVX1_35/Y BUFX4_23/Y gnd AOI21X1_59/C vdd OAI21X1
XNAND2X1_2 INVX1_19/A BUFX4_45/Y gnd OAI21X1_2/C vdd NAND2X1
XAOI21X1_7 INVX4_6/Y NOR2X1_9/B NOR2X1_9/Y gnd AOI21X1_7/Y vdd AOI21X1
XFILL_8_2_1 gnd vdd FILL
XINVX1_50 INVX1_50/A gnd INVX1_50/Y vdd INVX1
XFILL_0_1_1 gnd vdd FILL
XFILL_16_1_1 gnd vdd FILL
XNOR2X1_5 NOR2X1_5/A NOR2X1_9/B gnd NOR2X1_5/Y vdd NOR2X1
XBUFX2_14 INVX2_1/A gnd fifo_counter[4] vdd BUFX2
XDFFPOSX1_2 AOI21X1_41/B CLKBUF1_7/Y DFFPOSX1_2/D gnd vdd DFFPOSX1
XAOI21X1_15 OAI21X1_6/B NOR2X1_12/Y NOR2X1_18/Y gnd AOI21X1_15/Y vdd AOI21X1
XAOI21X1_26 rd_en INVX1_2/A AOI21X1_26/C gnd AOI21X1_26/Y vdd AOI21X1
XAOI21X1_37 NOR2X1_13/A BUFX4_2/Y BUFX4_23/Y gnd OAI21X1_71/C vdd AOI21X1
XOAI22X1_12 OAI22X1_12/A OAI22X1_12/B NAND2X1_71/Y BUFX4_34/Y gnd DFFSR_15/D vdd OAI22X1
XAOI21X1_48 BUFX4_41/Y INVX1_25/Y BUFX4_19/Y gnd OAI21X1_86/C vdd AOI21X1
XAOI21X1_59 BUFX4_26/Y AOI21X1_59/B AOI21X1_59/C gnd AOI21X1_59/Y vdd AOI21X1
XFILL_5_0_1 gnd vdd FILL
XDFFPOSX1_59 NAND2X1_78/A CLKBUF1_5/Y DFFPOSX1_59/D gnd vdd DFFPOSX1
XDFFPOSX1_37 INVX1_34/A CLKBUF1_5/Y OAI21X1_5/Y gnd vdd DFFPOSX1
XDFFPOSX1_26 NOR2X1_22/A CLKBUF1_12/Y AOI21X1_18/Y gnd vdd DFFPOSX1
XDFFPOSX1_48 NOR2X1_20/A CLKBUF1_9/Y AOI21X1_17/Y gnd vdd DFFPOSX1
XDFFPOSX1_15 INVX1_47/A CLKBUF1_1/Y MUX2X1_20/Y gnd vdd DFFPOSX1
XBUFX2_8 BUFX2_8/A gnd d_out[7] vdd BUFX2
XNOR2X1_70 NOR2X1_70/A NOR2X1_66/Y gnd NOR2X1_70/Y vdd NOR2X1
XAOI21X1_8 INVX4_7/Y NOR2X1_9/B NOR2X1_10/Y gnd AOI21X1_8/Y vdd AOI21X1
XNAND2X1_3 NOR2X1_40/A BUFX4_46/Y gnd OAI21X1_3/C vdd NAND2X1
XBUFX2_15 INVX1_1/Y gnd full vdd BUFX2
XINVX1_40 INVX1_40/A gnd INVX1_40/Y vdd INVX1
XNOR2X1_6 NOR2X1_6/A NOR2X1_9/B gnd NOR2X1_6/Y vdd NOR2X1
XDFFPOSX1_3 NOR2X1_41/A CLKBUF1_5/Y DFFPOSX1_3/D gnd vdd DFFPOSX1
XINVX1_51 INVX1_51/A gnd INVX1_51/Y vdd INVX1
XAOI21X1_27 INVX2_1/A NOR2X1_36/Y DFFSR_20/Q gnd AOI22X1_2/B vdd AOI21X1
XAOI21X1_38 OAI21X1_70/Y AOI21X1_38/B DFFSR_3/Q gnd OR2X2_1/B vdd AOI21X1
XAOI21X1_16 OAI21X1_7/B NOR2X1_12/Y NOR2X1_19/Y gnd AOI21X1_16/Y vdd AOI21X1
XAOI21X1_49 INVX8_2/A INVX1_26/Y BUFX4_18/Y gnd OAI21X1_91/C vdd AOI21X1
XOAI22X1_13 NOR2X1_55/Y OAI22X1_13/B OAI22X1_13/C NOR2X1_54/Y gnd OAI22X1_13/Y vdd
+ OAI22X1
XOAI21X1_90 BUFX4_39/Y NOR2X1_23/A INVX8_3/A gnd OAI22X1_3/B vdd OAI21X1
XDFFPOSX1_16 INVX1_53/A CLKBUF1_10/Y MUX2X1_21/Y gnd vdd DFFPOSX1
XDFFPOSX1_27 NOR2X1_23/A CLKBUF1_12/Y AOI21X1_19/Y gnd vdd DFFPOSX1
XDFFPOSX1_38 INVX1_40/A CLKBUF1_6/Y OAI21X1_6/Y gnd vdd DFFPOSX1
XDFFPOSX1_49 INVX1_10/A CLKBUF1_10/Y MUX2X1_1/Y gnd vdd DFFPOSX1
XFILL_14_2_0 gnd vdd FILL
XFILL_3_1_0 gnd vdd FILL
XNOR2X1_60 NOR2X1_60/A NOR2X1_58/Y gnd NOR2X1_60/Y vdd NOR2X1
XFILL_11_0_0 gnd vdd FILL
XNOR2X1_71 NOR2X1_71/A NOR2X1_66/Y gnd NOR2X1_71/Y vdd NOR2X1
XBUFX2_9 INVX1_2/Y gnd empty vdd BUFX2
XNAND2X1_4 INVX1_28/A BUFX4_44/Y gnd OAI21X1_4/C vdd NAND2X1
XAOI21X1_9 INVX4_8/Y NOR2X1_9/B AOI21X1_9/C gnd AOI21X1_9/Y vdd AOI21X1
XINVX1_41 INVX1_41/A gnd INVX1_41/Y vdd INVX1
XINVX1_52 INVX1_52/A gnd INVX1_52/Y vdd INVX1
XNOR2X1_7 NOR2X1_7/A NOR2X1_9/B gnd NOR2X1_7/Y vdd NOR2X1
XDFFPOSX1_4 NAND2X1_93/A CLKBUF1_11/Y DFFPOSX1_4/D gnd vdd DFFPOSX1
XINVX1_30 INVX1_30/A gnd INVX1_30/Y vdd INVX1
XAOI21X1_39 BUFX4_34/Y OR2X2_1/Y AOI21X1_32/Y gnd DFFSR_9/D vdd AOI21X1
XAOI21X1_17 OAI21X1_8/A NOR2X1_12/Y NOR2X1_20/Y gnd AOI21X1_17/Y vdd AOI21X1
XAOI21X1_28 BUFX4_27/Y NOR2X1_67/A AOI21X1_28/C gnd AOI21X1_28/Y vdd AOI21X1
XOAI22X1_14 OAI22X1_14/A OAI22X1_14/B NAND2X1_72/Y BUFX4_36/Y gnd DFFSR_16/D vdd OAI22X1
XFILL_8_0_0 gnd vdd FILL
XOAI21X1_80 BUFX4_24/Y NOR2X1_14/A BUFX4_3/Y gnd OAI22X1_1/C vdd OAI21X1
XOAI21X1_91 BUFX4_41/Y OAI21X1_91/B OAI21X1_91/C gnd OAI21X1_91/Y vdd OAI21X1
XDFFPOSX1_39 INVX1_46/A CLKBUF1_3/Y OAI21X1_7/Y gnd vdd DFFPOSX1
XDFFPOSX1_28 INVX1_31/A CLKBUF1_1/Y MUX2X1_9/Y gnd vdd DFFPOSX1
XDFFPOSX1_17 NOR2X1_59/A CLKBUF1_7/Y AOI21X1_85/Y gnd vdd DFFPOSX1
XFILL_14_2_1 gnd vdd FILL
XFILL_3_1_1 gnd vdd FILL
XNOR2X1_72 NOR2X1_72/A NOR2X1_66/Y gnd NOR2X1_72/Y vdd NOR2X1
XNOR2X1_50 BUFX4_38/Y NOR2X1_9/A gnd OAI22X1_9/D vdd NOR2X1
XFILL_11_0_1 gnd vdd FILL
XNOR2X1_61 NOR2X1_61/A NOR2X1_58/Y gnd NOR2X1_61/Y vdd NOR2X1
XNAND2X1_5 INVX1_34/A BUFX4_46/Y gnd OAI21X1_5/C vdd NAND2X1
XDFFPOSX1_5 AOI21X1_58/B CLKBUF1_3/Y DFFPOSX1_5/D gnd vdd DFFPOSX1
XINVX1_42 INVX1_42/A gnd INVX1_42/Y vdd INVX1
XINVX1_31 INVX1_31/A gnd INVX1_31/Y vdd INVX1
XINVX1_20 INVX1_20/A gnd INVX1_20/Y vdd INVX1
XINVX1_53 INVX1_53/A gnd INVX1_53/Y vdd INVX1
XNOR2X1_8 NOR2X1_8/A NOR2X1_9/B gnd NOR2X1_8/Y vdd NOR2X1
XAOI21X1_29 BUFX4_30/Y AOI21X1_29/B AOI21X1_29/C gnd AOI21X1_29/Y vdd AOI21X1
XAOI21X1_18 INVX4_2/Y MUX2X1_9/S NOR2X1_22/Y gnd AOI21X1_18/Y vdd AOI21X1
XFILL_8_0_1 gnd vdd FILL
XOAI21X1_81 BUFX4_43/Y NOR2X1_22/A BUFX4_16/Y gnd OAI22X1_1/B vdd OAI21X1
XOAI21X1_70 BUFX4_1/Y INVX1_16/Y AOI21X1_36/Y gnd OAI21X1_70/Y vdd OAI21X1
XOAI21X1_92 BUFX4_42/Y NAND2X1_38/A BUFX4_19/Y gnd OAI21X1_92/Y vdd OAI21X1
XDFFPOSX1_18 NOR2X1_60/A CLKBUF1_6/Y AOI21X1_86/Y gnd vdd DFFPOSX1
XDFFPOSX1_29 INVX1_37/A CLKBUF1_3/Y MUX2X1_10/Y gnd vdd DFFPOSX1
XNAND2X1_6 INVX1_40/A BUFX4_45/Y gnd OAI21X1_6/C vdd NAND2X1
XNOR2X1_51 NOR2X1_51/A BUFX4_21/Y gnd OAI22X1_9/A vdd NOR2X1
XNOR2X1_40 NOR2X1_40/A BUFX4_25/Y gnd NOR2X1_40/Y vdd NOR2X1
XNOR2X1_62 NOR2X1_62/A NOR2X1_58/Y gnd NOR2X1_62/Y vdd NOR2X1
XNOR2X1_73 NOR2X1_73/A NOR2X1_66/Y gnd NOR2X1_73/Y vdd NOR2X1
XDFFPOSX1_6 NAND2X1_95/A CLKBUF1_6/Y DFFPOSX1_6/D gnd vdd DFFPOSX1
XINVX1_21 INVX1_21/A gnd INVX1_21/Y vdd INVX1
XINVX1_43 INVX1_43/A gnd INVX1_43/Y vdd INVX1
XINVX1_32 INVX1_32/A gnd INVX1_32/Y vdd INVX1
XINVX1_10 INVX1_10/A gnd MUX2X1_1/B vdd INVX1
XINVX1_54 INVX1_54/A gnd INVX1_54/Y vdd INVX1
XNOR2X1_9 NOR2X1_9/A NOR2X1_9/B gnd NOR2X1_9/Y vdd NOR2X1
XAOI21X1_19 INVX4_3/Y MUX2X1_9/S NOR2X1_23/Y gnd AOI21X1_19/Y vdd AOI21X1
XOAI21X1_60 XNOR2X1_1/A NAND2X1_64/Y AOI22X1_2/A gnd AOI22X1_2/C vdd OAI21X1
XOAI21X1_71 BUFX4_2/Y INVX1_17/Y OAI21X1_71/C gnd AOI21X1_38/B vdd OAI21X1
XOAI21X1_82 OAI22X1_1/Y DFFSR_3/Q BUFX4_35/Y gnd OAI22X1_2/A vdd OAI21X1
XOAI21X1_93 NOR2X1_45/Y OAI21X1_92/Y OAI21X1_91/Y gnd OAI21X1_93/Y vdd OAI21X1
XFILL_1_2_0 gnd vdd FILL
XFILL_17_2_0 gnd vdd FILL
XDFFPOSX1_19 INVX1_25/A CLKBUF1_9/Y MUX2X1_14/Y gnd vdd DFFPOSX1
XFILL_14_0_0 gnd vdd FILL
XFILL_6_1_0 gnd vdd FILL
XNOR2X1_63 NOR2X1_63/A NOR2X1_58/Y gnd NOR2X1_63/Y vdd NOR2X1
XNOR2X1_30 XNOR2X1_5/A BUFX4_7/Y gnd NOR2X1_30/Y vdd NOR2X1
XNAND2X1_7 INVX1_46/A BUFX4_47/Y gnd NAND2X1_7/Y vdd NAND2X1
XNOR2X1_41 NOR2X1_41/A BUFX4_25/Y gnd NOR2X1_41/Y vdd NOR2X1
XNOR2X1_74 NOR2X1_74/A NOR2X1_66/Y gnd NOR2X1_74/Y vdd NOR2X1
XNOR2X1_52 BUFX4_43/Y NOR2X1_52/B gnd NOR2X1_52/Y vdd NOR2X1
XINVX1_22 INVX1_22/A gnd INVX1_22/Y vdd INVX1
XINVX1_33 INVX1_33/A gnd MUX2X1_4/B vdd INVX1
XINVX1_11 INVX1_11/A gnd INVX1_11/Y vdd INVX1
XINVX1_55 INVX1_55/A gnd INVX1_55/Y vdd INVX1
XINVX1_44 INVX1_44/A gnd INVX1_44/Y vdd INVX1
XDFFPOSX1_7 AOI21X1_72/B CLKBUF1_5/Y DFFPOSX1_7/D gnd vdd DFFPOSX1
XOAI21X1_50 NOR2X1_36/B INVX2_1/A rd_en gnd XNOR2X1_5/A vdd OAI21X1
XOAI21X1_61 OAI21X1_61/A AOI21X1_26/C OAI21X1_61/C gnd AOI22X1_3/C vdd OAI21X1
XOAI21X1_83 BUFX4_39/Y NOR2X1_76/A OAI21X1_83/C gnd OAI21X1_85/C vdd OAI21X1
XOAI21X1_72 BUFX4_26/Y INVX1_18/Y BUFX4_24/Y gnd AOI21X1_40/C vdd OAI21X1
XOAI21X1_94 OAI21X1_93/Y BUFX4_30/Y BUFX4_37/Y gnd OAI22X1_4/A vdd OAI21X1
XFILL_1_2_1 gnd vdd FILL
XFILL_17_2_1 gnd vdd FILL
XDFFSR_20 DFFSR_20/Q CLKBUF1_2/Y DFFSR_5/R vdd DFFSR_20/D gnd vdd DFFSR
XFILL_14_0_1 gnd vdd FILL
XFILL_6_1_1 gnd vdd FILL
XNOR2X1_75 NOR2X1_75/A NOR2X1_3/B gnd MUX2X1_19/S vdd NOR2X1
XNOR2X1_31 BUFX4_23/Y BUFX4_2/Y gnd INVX1_5/A vdd NOR2X1
XNOR2X1_42 BUFX4_38/Y NOR2X1_6/A gnd OAI22X1_3/D vdd NOR2X1
XNOR2X1_53 NOR2X1_53/A BUFX4_25/Y gnd NOR2X1_53/Y vdd NOR2X1
XNOR2X1_20 NOR2X1_20/A NOR2X1_12/Y gnd NOR2X1_20/Y vdd NOR2X1
XNOR2X1_64 NOR2X1_64/A NOR2X1_58/Y gnd NOR2X1_64/Y vdd NOR2X1
XNAND2X1_8 INVX1_52/A BUFX4_47/Y gnd NAND2X1_8/Y vdd NAND2X1
XINVX1_23 INVX1_23/A gnd INVX1_23/Y vdd INVX1
XINVX1_45 INVX1_45/A gnd INVX1_45/Y vdd INVX1
XDFFPOSX1_8 DFFPOSX1_8/Q CLKBUF1_11/Y DFFPOSX1_8/D gnd vdd DFFPOSX1
XINVX1_34 INVX1_34/A gnd INVX1_34/Y vdd INVX1
XINVX1_12 INVX1_12/A gnd INVX1_12/Y vdd INVX1
XINVX1_56 INVX1_56/A gnd INVX1_56/Y vdd INVX1
XOAI21X1_40 OAI21X1_8/A NAND3X1_4/Y OAI21X1_40/C gnd OAI21X1_40/Y vdd OAI21X1
XOAI21X1_51 XNOR2X1_1/A INVX1_5/Y DFFSR_3/Q gnd OAI21X1_51/Y vdd OAI21X1
XOAI21X1_73 BUFX4_31/Y INVX1_19/Y BUFX4_39/Y gnd AOI21X1_41/C vdd OAI21X1
XOAI21X1_84 INVX8_2/A NOR2X1_1/A BUFX4_18/Y gnd OAI21X1_85/B vdd OAI21X1
XOAI21X1_62 BUFX4_27/Y MUX2X1_1/B BUFX4_22/Y gnd AOI21X1_28/C vdd OAI21X1
XOAI21X1_95 BUFX4_27/Y MUX2X1_3/B BUFX4_22/Y gnd AOI21X1_50/C vdd OAI21X1
XDFFSR_21 INVX2_1/A CLKBUF1_2/Y DFFSR_1/R vdd DFFSR_21/D gnd vdd DFFSR
XDFFSR_10 BUFX2_2/A CLKBUF1_8/Y DFFSR_9/R vdd DFFSR_10/D gnd vdd DFFSR
XFILL_18_1 gnd vdd FILL
XNAND3X1_10 wr_en XOR2X1_1/Y INVX1_1/A gnd INVX1_6/A vdd NAND3X1
XNOR2X1_32 INVX1_4/A INVX2_3/Y gnd NOR2X1_32/Y vdd NOR2X1
XNOR2X1_21 NOR2X1_21/A NOR2X1_3/B gnd MUX2X1_9/S vdd NOR2X1
XNOR2X1_10 NOR2X1_10/A NOR2X1_9/B gnd NOR2X1_10/Y vdd NOR2X1
XNOR2X1_54 BUFX4_42/Y NOR2X1_11/A gnd NOR2X1_54/Y vdd NOR2X1
XNOR2X1_76 NOR2X1_76/A MUX2X1_19/S gnd NOR2X1_76/Y vdd NOR2X1
XNOR2X1_65 NOR2X1_65/A NOR2X1_58/Y gnd NOR2X1_65/Y vdd NOR2X1
XNOR2X1_43 NOR2X1_43/A BUFX4_24/Y gnd NOR2X1_43/Y vdd NOR2X1
XNAND2X1_9 NOR2X1_57/Y NOR2X1_2/Y gnd NOR2X1_3/A vdd NAND2X1
XINVX1_13 INVX1_13/A gnd INVX1_13/Y vdd INVX1
XINVX1_35 INVX1_35/A gnd INVX1_35/Y vdd INVX1
XINVX1_46 INVX1_46/A gnd INVX1_46/Y vdd INVX1
XINVX1_24 INVX1_24/A gnd INVX1_24/Y vdd INVX1
XDFFPOSX1_9 INVX1_12/A CLKBUF1_10/Y MUX2X1_15/Y gnd vdd DFFPOSX1
XFILL_12_1_0 gnd vdd FILL
XFILL_4_2_0 gnd vdd FILL
XOAI21X1_30 OAI21X1_6/B NAND3X1_3/Y NAND2X1_33/Y gnd OAI21X1_30/Y vdd OAI21X1
XOAI21X1_52 MUX2X1_12/Y BUFX4_9/Y NAND2X1_57/Y gnd DFFSR_4/D vdd OAI21X1
XOAI21X1_41 NAND3X1_7/Y OAI21X1_9/A OAI21X1_41/C gnd OAI21X1_41/Y vdd OAI21X1
XOAI21X1_63 BUFX4_30/Y INVX1_11/Y BUFX4_41/Y gnd AOI21X1_29/C vdd OAI21X1
XOAI21X1_96 BUFX4_29/Y INVX1_28/Y BUFX4_43/Y gnd OAI21X1_96/Y vdd OAI21X1
XOAI21X1_85 NOR2X1_40/Y OAI21X1_85/B OAI21X1_85/C gnd MUX2X1_13/B vdd OAI21X1
XOAI21X1_74 AOI21X1_40/Y OAI21X1_74/B BUFX4_19/Y gnd OAI21X1_74/Y vdd OAI21X1
XDFFSR_11 BUFX2_3/A CLKBUF1_6/Y DFFSR_4/R vdd DFFSR_11/D gnd vdd DFFSR
XFILL_1_0_0 gnd vdd FILL
XFILL_17_0_0 gnd vdd FILL
XFILL_9_1_0 gnd vdd FILL
XNOR2X1_33 DFFSR_6/Q INVX1_4/Y gnd NOR2X1_33/Y vdd NOR2X1
XNAND3X1_11 rd_en XNOR2X1_7/Y INVX1_2/A gnd OAI21X1_56/C vdd NAND3X1
XNOR2X1_66 NOR2X1_66/A NOR2X1_3/B gnd NOR2X1_66/Y vdd NOR2X1
XNOR2X1_77 NOR2X1_77/A NOR2X1_3/B gnd NOR2X1_77/Y vdd NOR2X1
XNOR2X1_11 NOR2X1_11/A NOR2X1_9/B gnd AOI21X1_9/C vdd NOR2X1
XNOR2X1_44 DFFSR_3/Q OAI22X1_3/Y gnd OAI22X1_4/B vdd NOR2X1
XNOR2X1_22 NOR2X1_22/A MUX2X1_9/S gnd NOR2X1_22/Y vdd NOR2X1
XNOR2X1_55 NOR2X1_55/A BUFX4_24/Y gnd NOR2X1_55/Y vdd NOR2X1
XINVX1_36 INVX1_36/A gnd INVX1_36/Y vdd INVX1
XINVX1_25 INVX1_25/A gnd INVX1_25/Y vdd INVX1
XINVX1_14 INVX1_14/A gnd INVX1_14/Y vdd INVX1
XINVX1_47 INVX1_47/A gnd INVX1_47/Y vdd INVX1
XFILL_12_1_1 gnd vdd FILL
XFILL_4_2_1 gnd vdd FILL
XOAI21X1_53 NOR2X1_32/Y NOR2X1_33/Y BUFX4_11/Y gnd OAI21X1_53/Y vdd OAI21X1
XOAI21X1_42 NAND3X1_7/Y OAI21X1_2/B NAND2X1_45/Y gnd OAI21X1_42/Y vdd OAI21X1
XOAI21X1_20 OAI21X1_4/B NAND3X1_2/Y OAI21X1_20/C gnd OAI21X1_20/Y vdd OAI21X1
XOAI21X1_64 AOI21X1_28/Y AOI21X1_29/Y BUFX4_18/Y gnd OAI21X1_64/Y vdd OAI21X1
XOAI21X1_86 BUFX4_42/Y NAND2X1_78/A OAI21X1_86/C gnd OAI21X1_86/Y vdd OAI21X1
XOAI21X1_75 BUFX4_33/Y INVX1_20/Y BUFX4_25/Y gnd AOI21X1_42/C vdd OAI21X1
XOAI21X1_97 OAI21X1_97/A OAI21X1_97/B BUFX4_16/Y gnd NAND2X1_68/A vdd OAI21X1
XOAI21X1_31 OAI21X1_7/B NAND3X1_3/Y NAND2X1_34/Y gnd OAI21X1_31/Y vdd OAI21X1
XDFFSR_12 BUFX2_4/A CLKBUF1_6/Y DFFSR_4/R vdd DFFSR_12/D gnd vdd DFFSR
XCLKBUF1_10 clk gnd CLKBUF1_10/Y vdd CLKBUF1
XFILL_1_0_1 gnd vdd FILL
XFILL_17_0_1 gnd vdd FILL
XFILL_9_1_1 gnd vdd FILL
XNOR2X1_12 NOR2X1_12/A NOR2X1_3/B gnd NOR2X1_12/Y vdd NOR2X1
XNAND3X1_12 AND2X2_3/Y XNOR2X1_5/A BUFX4_8/Y gnd AOI22X1_1/D vdd NAND3X1
XNOR2X1_56 INVX1_3/A DFFSR_7/Q gnd NOR2X1_56/Y vdd NOR2X1
XNOR2X1_34 INVX1_3/A INVX2_2/Y gnd NOR2X1_34/Y vdd NOR2X1
XNOR2X1_78 NOR2X1_78/A NOR2X1_3/B gnd MUX2X1_5/S vdd NOR2X1
XNOR2X1_45 NOR2X1_45/A BUFX4_25/Y gnd NOR2X1_45/Y vdd NOR2X1
XNOR2X1_67 NOR2X1_67/A NOR2X1_66/Y gnd NOR2X1_67/Y vdd NOR2X1
XNOR2X1_23 NOR2X1_23/A MUX2X1_9/S gnd NOR2X1_23/Y vdd NOR2X1
XINVX1_37 INVX1_37/A gnd INVX1_37/Y vdd INVX1
XINVX1_15 INVX1_15/A gnd INVX1_15/Y vdd INVX1
XINVX1_26 INVX1_26/A gnd INVX1_26/Y vdd INVX1
XINVX1_48 INVX1_48/A gnd INVX1_48/Y vdd INVX1
XOAI21X1_54 INVX2_3/Y BUFX4_11/Y OAI21X1_53/Y gnd DFFSR_6/D vdd OAI21X1
XOAI21X1_76 BUFX4_32/Y INVX1_21/Y INVX8_2/A gnd OAI21X1_76/Y vdd OAI21X1
XOAI21X1_32 OAI21X1_8/A NAND3X1_3/Y NAND2X1_35/Y gnd OAI21X1_32/Y vdd OAI21X1
XOAI21X1_21 MUX2X1_26/A NAND3X1_2/Y NAND2X1_24/Y gnd OAI21X1_21/Y vdd OAI21X1
XOAI21X1_10 OAI21X1_2/B NAND3X1_1/Y NAND2X1_13/Y gnd OAI21X1_10/Y vdd OAI21X1
XOAI21X1_43 NAND3X1_7/Y MUX2X1_24/A NAND2X1_46/Y gnd OAI21X1_43/Y vdd OAI21X1
XOAI21X1_87 BUFX4_43/Y NOR2X1_69/A BUFX4_16/Y gnd OAI21X1_88/B vdd OAI21X1
XOAI21X1_98 BUFX4_26/Y INVX1_29/Y BUFX4_24/Y gnd OAI21X1_98/Y vdd OAI21X1
XOAI21X1_65 BUFX4_29/Y INVX1_12/Y BUFX4_20/Y gnd AOI21X1_30/C vdd OAI21X1
XDFFSR_13 BUFX2_5/A CLKBUF1_6/Y DFFSR_9/R vdd DFFSR_13/D gnd vdd DFFSR
XCLKBUF1_11 clk gnd CLKBUF1_11/Y vdd CLKBUF1
XFILL_10_2_0 gnd vdd FILL
XNOR2X1_35 NOR2X1_3/B XNOR2X1_5/A gnd NOR2X1_35/Y vdd NOR2X1
XNOR2X1_57 DFFSR_6/Q INVX1_4/A gnd NOR2X1_57/Y vdd NOR2X1
XNAND3X1_13 DFFSR_20/Q AOI21X1_26/Y BUFX4_8/Y gnd AOI22X1_3/B vdd NAND3X1
XNOR2X1_24 NOR2X1_24/A MUX2X1_9/S gnd NOR2X1_24/Y vdd NOR2X1
XNOR2X1_46 INVX8_2/A NOR2X1_46/B gnd OAI22X1_5/D vdd NOR2X1
XNOR2X1_13 NOR2X1_13/A NOR2X1_12/Y gnd NOR2X1_13/Y vdd NOR2X1
XNOR2X1_68 NOR2X1_68/A NOR2X1_66/Y gnd NOR2X1_68/Y vdd NOR2X1
XFILL_16_1 gnd vdd FILL
XDFFSR_1 DFFSR_1/Q CLKBUF1_2/Y DFFSR_1/R vdd DFFSR_1/D gnd vdd DFFSR
XINVX1_38 INVX1_38/A gnd INVX1_38/Y vdd INVX1
XINVX1_49 INVX1_49/A gnd INVX1_49/Y vdd INVX1
XINVX1_16 INVX1_16/A gnd INVX1_16/Y vdd INVX1
XINVX1_27 INVX1_27/A gnd MUX2X1_3/B vdd INVX1
XMUX2X1_20 INVX4_7/Y INVX1_47/Y MUX2X1_19/S gnd MUX2X1_20/Y vdd MUX2X1
XNAND2X1_90 AOI21X1_29/B NAND3X1_15/Y gnd NAND2X1_90/Y vdd NAND2X1
XFILL_7_2_0 gnd vdd FILL
XFILL_15_1_0 gnd vdd FILL
XOAI21X1_55 XNOR2X1_4/A INVX2_2/Y INVX1_3/A gnd NAND2X1_59/B vdd OAI21X1
XOAI21X1_44 NAND3X1_7/Y OAI21X1_4/B NAND2X1_47/Y gnd OAI21X1_44/Y vdd OAI21X1
XOAI21X1_66 BUFX4_30/Y INVX1_13/Y BUFX4_42/Y gnd OAI21X1_66/Y vdd OAI21X1
XOAI21X1_11 MUX2X1_24/A NAND3X1_1/Y NAND2X1_14/Y gnd OAI21X1_11/Y vdd OAI21X1
XOAI21X1_88 NOR2X1_41/Y OAI21X1_88/B OAI21X1_86/Y gnd MUX2X1_13/A vdd OAI21X1
XOAI21X1_99 BUFX4_33/Y INVX1_30/Y BUFX4_38/Y gnd OAI21X1_99/Y vdd OAI21X1
XOAI21X1_33 OAI21X1_9/A NAND3X1_4/Y NAND2X1_36/Y gnd OAI21X1_33/Y vdd OAI21X1
XOAI21X1_77 AOI21X1_42/Y OAI21X1_77/B BUFX4_6/Y gnd OAI21X1_77/Y vdd OAI21X1
XOAI21X1_22 OAI21X1_6/B NAND3X1_2/Y OAI21X1_22/C gnd OAI21X1_22/Y vdd OAI21X1
XFILL_4_0_0 gnd vdd FILL
XDFFSR_14 BUFX2_6/A CLKBUF1_8/Y DFFSR_9/R vdd DFFSR_14/D gnd vdd DFFSR
XCLKBUF1_12 clk gnd CLKBUF1_12/Y vdd CLKBUF1
XFILL_4_1 gnd vdd FILL
XFILL_10_2_1 gnd vdd FILL
XNOR2X1_58 NOR2X1_58/A NOR2X1_3/B gnd NOR2X1_58/Y vdd NOR2X1
XNOR2X1_36 INVX1_8/Y NOR2X1_36/B gnd NOR2X1_36/Y vdd NOR2X1
XNAND3X1_14 NOR2X1_56/Y NOR2X1_57/Y BUFX4_7/Y gnd NAND3X1_14/Y vdd NAND3X1
XNOR2X1_47 NOR2X1_47/A BUFX4_21/Y gnd OAI22X1_5/A vdd NOR2X1
XNOR2X1_25 NOR2X1_25/A MUX2X1_9/S gnd NOR2X1_25/Y vdd NOR2X1
XNOR2X1_14 NOR2X1_14/A NOR2X1_12/Y gnd NOR2X1_14/Y vdd NOR2X1
XNOR2X1_69 NOR2X1_69/A NOR2X1_66/Y gnd NOR2X1_69/Y vdd NOR2X1
XDFFSR_2 DFFSR_2/Q CLKBUF1_3/Y DFFSR_1/R vdd DFFSR_2/D gnd vdd DFFSR
XMUX2X1_10 INVX4_5/Y INVX1_37/Y MUX2X1_9/S gnd MUX2X1_10/Y vdd MUX2X1
XMUX2X1_21 INVX4_8/Y INVX1_53/Y MUX2X1_19/S gnd MUX2X1_21/Y vdd MUX2X1
XINVX1_39 INVX1_39/A gnd INVX1_39/Y vdd INVX1
XINVX1_17 INVX1_17/A gnd INVX1_17/Y vdd INVX1
XINVX1_28 INVX1_28/A gnd INVX1_28/Y vdd INVX1
XFILL_7_2_1 gnd vdd FILL
XNAND2X1_80 AOI21X1_52/B NAND3X1_14/Y gnd NAND2X1_80/Y vdd NAND2X1
XNAND2X1_91 AOI21X1_41/B NAND3X1_15/Y gnd NAND2X1_91/Y vdd NAND2X1
XFILL_15_1_1 gnd vdd FILL
XOAI21X1_34 OAI21X1_2/B NAND3X1_4/Y NAND2X1_37/Y gnd OAI21X1_34/Y vdd OAI21X1
XOAI21X1_45 NAND3X1_7/Y MUX2X1_26/A OAI21X1_45/C gnd OAI21X1_45/Y vdd OAI21X1
XOAI21X1_12 OAI21X1_4/B NAND3X1_1/Y NAND2X1_15/Y gnd OAI21X1_12/Y vdd OAI21X1
XOAI21X1_23 OAI21X1_7/B NAND3X1_2/Y OAI21X1_23/C gnd OAI21X1_23/Y vdd OAI21X1
XOAI21X1_56 AND2X2_2/Y INVX1_7/Y OAI21X1_56/C gnd AOI21X1_24/B vdd OAI21X1
XOAI21X1_78 BUFX4_4/Y INVX1_22/Y AOI21X1_44/Y gnd AOI21X1_46/A vdd OAI21X1
XOAI21X1_67 AOI21X1_30/Y AOI21X1_31/Y BUFX4_6/Y gnd OAI21X1_67/Y vdd OAI21X1
XOAI21X1_89 BUFX4_24/Y NOR2X1_15/A BUFX4_3/Y gnd OAI22X1_3/C vdd OAI21X1
XFILL_4_0_1 gnd vdd FILL
XDFFSR_15 BUFX2_7/A CLKBUF1_8/Y DFFSR_9/R vdd DFFSR_15/D gnd vdd DFFSR
XNOR2X1_37 INVX2_1/Y NOR2X1_35/Y gnd AOI22X1_3/D vdd NOR2X1
XNOR2X1_26 INVX1_7/A DFFSR_17/Q gnd NAND3X1_5/B vdd NOR2X1
XNAND3X1_15 NOR2X1_29/Y NOR2X1_56/Y BUFX4_9/Y gnd NAND3X1_15/Y vdd NAND3X1
XNOR2X1_15 NOR2X1_15/A NOR2X1_12/Y gnd NOR2X1_15/Y vdd NOR2X1
XNOR2X1_48 BUFX4_39/Y NOR2X1_48/B gnd NOR2X1_48/Y vdd NOR2X1
XNOR2X1_59 NOR2X1_59/A NOR2X1_58/Y gnd NOR2X1_59/Y vdd NOR2X1
XDFFSR_3 DFFSR_3/Q CLKBUF1_2/Y DFFSR_1/R vdd DFFSR_3/D gnd vdd DFFSR
XMUX2X1_22 OAI21X1_9/A INVX1_13/Y NOR2X1_77/Y gnd MUX2X1_22/Y vdd MUX2X1
XMUX2X1_11 INVX4_7/Y INVX1_49/Y MUX2X1_9/S gnd MUX2X1_11/Y vdd MUX2X1
XNAND2X1_70 NAND2X1_70/A NAND2X1_70/B gnd OAI22X1_10/C vdd NAND2X1
XNAND2X1_81 d_in[4] BUFX4_10/Y gnd MUX2X1_26/A vdd NAND2X1
XINVX1_18 INVX1_18/A gnd INVX1_18/Y vdd INVX1
XNAND2X1_92 NOR2X1_41/A NAND3X1_15/Y gnd NAND2X1_92/Y vdd NAND2X1
XINVX1_29 INVX1_29/A gnd INVX1_29/Y vdd INVX1
XOAI21X1_57 OAI21X1_57/A NOR2X1_35/Y OAI21X1_57/C gnd DFFSR_18/D vdd OAI21X1
XOAI21X1_24 OAI21X1_8/A NAND3X1_2/Y NAND2X1_27/Y gnd OAI21X1_24/Y vdd OAI21X1
XOAI21X1_13 MUX2X1_26/A NAND3X1_1/Y NAND2X1_16/Y gnd OAI21X1_13/Y vdd OAI21X1
XOAI21X1_79 BUFX4_4/Y INVX1_23/Y AOI21X1_45/Y gnd AOI21X1_46/B vdd OAI21X1
XOAI21X1_35 MUX2X1_24/A NAND3X1_4/Y OAI21X1_35/C gnd OAI21X1_35/Y vdd OAI21X1
XOAI21X1_68 BUFX4_3/Y INVX1_14/Y AOI21X1_33/Y gnd OAI21X1_68/Y vdd OAI21X1
XOAI21X1_46 NAND3X1_7/Y OAI21X1_6/B OAI21X1_46/C gnd OAI21X1_46/Y vdd OAI21X1
XDFFSR_16 BUFX2_8/A CLKBUF1_8/Y DFFSR_9/R vdd DFFSR_16/D gnd vdd DFFSR
XFILL_13_2_0 gnd vdd FILL
XNOR2X1_27 DFFSR_20/Q INVX1_9/A gnd NAND3X1_5/C vdd NOR2X1
XNOR2X1_49 NOR2X1_49/A BUFX4_21/Y gnd OAI22X1_7/A vdd NOR2X1
XNOR2X1_16 NOR2X1_16/A NOR2X1_12/Y gnd NOR2X1_16/Y vdd NOR2X1
XNOR2X1_38 BUFX4_42/Y NOR2X1_5/A gnd OAI22X1_1/D vdd NOR2X1
XFILL_2_1_0 gnd vdd FILL
XMUX2X1_12 XNOR2X1_2/Y BUFX4_35/Y AND2X2_2/Y gnd MUX2X1_12/Y vdd MUX2X1
XMUX2X1_23 OAI21X1_2/B INVX1_21/Y NOR2X1_77/Y gnd MUX2X1_23/Y vdd MUX2X1
XFILL_10_0_0 gnd vdd FILL
XNAND2X1_60 INVX1_7/A NOR2X1_35/Y gnd OAI21X1_57/C vdd NAND2X1
XINVX1_19 INVX1_19/A gnd INVX1_19/Y vdd INVX1
XDFFSR_4 DFFSR_4/Q CLKBUF1_6/Y DFFSR_4/R vdd DFFSR_4/D gnd vdd DFFSR
XNAND2X1_93 NAND2X1_93/A NAND3X1_15/Y gnd NAND2X1_93/Y vdd NAND2X1
XNAND2X1_71 NAND2X1_71/A NAND2X1_71/B gnd NAND2X1_71/Y vdd NAND2X1
XNAND2X1_82 AOI21X1_59/B NAND3X1_14/Y gnd NAND2X1_82/Y vdd NAND2X1
XFILL_14_1 gnd vdd FILL
XFILL_7_0_0 gnd vdd FILL
XOAI21X1_58 XNOR2X1_5/A NAND2X1_61/Y NOR2X1_3/B gnd AOI22X1_1/A vdd OAI21X1
XOAI21X1_14 OAI21X1_6/B NAND3X1_1/Y OAI21X1_14/C gnd OAI21X1_14/Y vdd OAI21X1
XOAI21X1_69 BUFX4_1/Y INVX1_15/Y OAI21X1_69/C gnd AOI21X1_35/B vdd OAI21X1
XOAI21X1_25 OAI21X1_9/A NAND3X1_3/Y NAND2X1_28/Y gnd OAI21X1_25/Y vdd OAI21X1
XOAI21X1_47 NAND3X1_7/Y OAI21X1_7/B OAI21X1_47/C gnd OAI21X1_47/Y vdd OAI21X1
XOAI21X1_36 OAI21X1_4/B NAND3X1_4/Y OAI21X1_36/C gnd OAI21X1_36/Y vdd OAI21X1
XDFFPOSX1_120 NAND2X1_27/A CLKBUF1_4/Y OAI21X1_24/Y gnd vdd DFFPOSX1
XDFFSR_17 DFFSR_17/Q CLKBUF1_2/Y DFFSR_5/R vdd DFFSR_17/D gnd vdd DFFSR
XINVX1_1 INVX1_1/A gnd INVX1_1/Y vdd INVX1
XXNOR2X1_1 XNOR2X1_1/A BUFX4_38/Y gnd DFFSR_1/D vdd XNOR2X1
XFILL_13_2_1 gnd vdd FILL
XAND2X2_1 INVX1_1/A wr_en gnd BUFX4_7/A vdd AND2X2
XFILL_2_1 gnd vdd FILL
XNOR2X1_28 INVX1_3/Y INVX2_2/Y gnd NAND3X1_4/A vdd NOR2X1
XNOR2X1_17 NOR2X1_17/A NOR2X1_12/Y gnd NOR2X1_17/Y vdd NOR2X1
XFILL_10_0_1 gnd vdd FILL
XNOR2X1_39 NOR2X1_39/A BUFX4_25/Y gnd NOR2X1_39/Y vdd NOR2X1
XMUX2X1_13 MUX2X1_13/A MUX2X1_13/B BUFX4_33/Y gnd MUX2X1_13/Y vdd MUX2X1
XFILL_2_1_1 gnd vdd FILL
XMUX2X1_24 MUX2X1_24/A INVX1_24/Y NOR2X1_77/Y gnd MUX2X1_24/Y vdd MUX2X1
XDFFSR_5 INVX1_4/A CLKBUF1_2/Y DFFSR_5/R vdd DFFSR_5/D gnd vdd DFFSR
XNAND2X1_61 INVX1_9/A NAND3X1_5/B gnd NAND2X1_61/Y vdd NAND2X1
XNAND2X1_94 AOI21X1_58/B NAND3X1_15/Y gnd NAND2X1_94/Y vdd NAND2X1
XNAND2X1_83 d_in[5] BUFX4_8/Y gnd OAI21X1_6/B vdd NAND2X1
XNAND2X1_50 NOR2X1_53/A NAND3X1_7/Y gnd OAI21X1_47/C vdd NAND2X1
XNAND2X1_72 NAND2X1_72/A NAND2X1_72/B gnd NAND2X1_72/Y vdd NAND2X1
XOAI21X1_59 AND2X2_2/Y AOI21X1_26/C BUFX4_7/Y gnd AOI22X1_1/B vdd OAI21X1
XOAI21X1_26 OAI21X1_2/B NAND3X1_3/Y NAND2X1_29/Y gnd OAI21X1_26/Y vdd OAI21X1
XOAI21X1_15 OAI21X1_7/B NAND3X1_1/Y OAI21X1_15/C gnd OAI21X1_15/Y vdd OAI21X1
XOAI21X1_37 MUX2X1_26/A NAND3X1_4/Y OAI21X1_37/C gnd OAI21X1_37/Y vdd OAI21X1
XOAI21X1_48 NAND3X1_7/Y OAI21X1_8/A NAND2X1_52/Y gnd OAI21X1_48/Y vdd OAI21X1
XFILL_7_0_1 gnd vdd FILL
XDFFPOSX1_110 AOI21X1_69/A CLKBUF1_8/Y OAI21X1_30/Y gnd vdd DFFPOSX1
XDFFPOSX1_121 INVX1_17/A CLKBUF1_3/Y OAI21X1_9/Y gnd vdd DFFPOSX1
XDFFSR_18 INVX1_7/A CLKBUF1_2/Y DFFSR_5/R vdd DFFSR_18/D gnd vdd DFFSR
XXNOR2X1_2 XNOR2X1_2/A BUFX4_34/Y gnd XNOR2X1_2/Y vdd XNOR2X1
XINVX1_2 INVX1_2/A gnd INVX1_2/Y vdd INVX1
XAND2X2_2 INVX1_2/A rd_en gnd AND2X2_2/Y vdd AND2X2
XFILL_2_2 gnd vdd FILL
XNOR2X1_29 INVX2_3/Y INVX1_4/Y gnd NOR2X1_29/Y vdd NOR2X1
XNOR2X1_18 NOR2X1_18/A NOR2X1_12/Y gnd NOR2X1_18/Y vdd NOR2X1
XDFFSR_6 DFFSR_6/Q CLKBUF1_2/Y DFFSR_5/R vdd DFFSR_6/D gnd vdd DFFSR
XNAND2X1_95 NAND2X1_95/A NAND3X1_15/Y gnd NAND2X1_95/Y vdd NAND2X1
XNAND2X1_62 INVX1_9/A AND2X2_3/Y gnd AOI21X1_26/C vdd NAND2X1
XNAND2X1_51 d_in[7] BUFX4_7/Y gnd OAI21X1_8/A vdd NAND2X1
XNAND2X1_84 AOI21X1_66/B NAND3X1_14/Y gnd NAND2X1_84/Y vdd NAND2X1
XMUX2X1_25 OAI21X1_4/B INVX1_30/Y NOR2X1_77/Y gnd MUX2X1_25/Y vdd MUX2X1
XMUX2X1_14 MUX2X1_24/A INVX1_25/Y NOR2X1_58/Y gnd MUX2X1_14/Y vdd MUX2X1
XNAND2X1_40 NAND2X1_40/A NAND3X1_4/Y gnd OAI21X1_37/C vdd NAND2X1
XNAND2X1_73 d_in[0] BUFX4_10/Y gnd OAI21X1_9/A vdd NAND2X1
XOAI21X1_49 NOR2X1_36/B INVX2_1/Y wr_en gnd NOR2X1_3/B vdd OAI21X1
XOAI21X1_38 OAI21X1_6/B NAND3X1_4/Y OAI21X1_38/C gnd OAI21X1_38/Y vdd OAI21X1
XOAI21X1_16 OAI21X1_8/A NAND3X1_1/Y OAI21X1_16/C gnd OAI21X1_16/Y vdd OAI21X1
XOAI21X1_27 MUX2X1_24/A NAND3X1_3/Y NAND2X1_30/Y gnd OAI21X1_27/Y vdd OAI21X1
XDFFPOSX1_100 INVX1_30/A CLKBUF1_5/Y MUX2X1_25/Y gnd vdd DFFPOSX1
XDFFPOSX1_122 NOR2X1_39/A CLKBUF1_5/Y OAI21X1_10/Y gnd vdd DFFPOSX1
XDFFPOSX1_111 NAND2X1_34/A CLKBUF1_7/Y OAI21X1_31/Y gnd vdd DFFPOSX1
XFILL_0_2_0 gnd vdd FILL
XFILL_16_2_0 gnd vdd FILL
XDFFSR_19 INVX1_9/A CLKBUF1_2/Y DFFSR_1/R vdd DFFSR_19/D gnd vdd DFFSR
XXNOR2X1_3 NOR2X1_3/B INVX1_4/A gnd DFFSR_5/D vdd XNOR2X1
XOR2X2_1 OR2X2_1/A OR2X2_1/B gnd OR2X2_1/Y vdd OR2X2
XINVX1_3 INVX1_3/A gnd INVX1_3/Y vdd INVX1
XFILL_13_0_0 gnd vdd FILL
XFILL_5_1_0 gnd vdd FILL
XAND2X2_3 INVX1_7/A DFFSR_17/Q gnd AND2X2_3/Y vdd AND2X2
XNOR2X1_19 NOR2X1_19/A NOR2X1_12/Y gnd NOR2X1_19/Y vdd NOR2X1
XDFFSR_7 DFFSR_7/Q CLKBUF1_3/Y DFFSR_4/R vdd DFFSR_7/D gnd vdd DFFSR
XMUX2X1_26 MUX2X1_26/A INVX1_36/Y NOR2X1_77/Y gnd MUX2X1_26/Y vdd MUX2X1
XMUX2X1_15 INVX4_1/Y INVX1_12/Y MUX2X1_19/S gnd MUX2X1_15/Y vdd MUX2X1
XNAND2X1_63 AOI21X1_26/Y BUFX4_8/Y gnd AOI22X1_2/A vdd NAND2X1
XNAND2X1_85 d_in[6] BUFX4_8/Y gnd OAI21X1_7/B vdd NAND2X1
XNAND2X1_41 INVX1_43/A NAND3X1_4/Y gnd OAI21X1_38/C vdd NAND2X1
XNAND2X1_96 AOI21X1_72/B NAND3X1_15/Y gnd NAND2X1_96/Y vdd NAND2X1
XNAND2X1_30 INVX1_26/A NAND3X1_3/Y gnd NAND2X1_30/Y vdd NAND2X1
XNAND2X1_52 INVX1_56/A NAND3X1_7/Y gnd NAND2X1_52/Y vdd NAND2X1
XNAND2X1_74 AOI21X1_30/B NAND3X1_14/Y gnd NAND2X1_74/Y vdd NAND2X1
XOAI22X1_1 NOR2X1_39/Y OAI22X1_1/B OAI22X1_1/C OAI22X1_1/D gnd OAI22X1_1/Y vdd OAI22X1
XOAI21X1_39 OAI21X1_7/B NAND3X1_4/Y OAI21X1_39/C gnd OAI21X1_39/Y vdd OAI21X1
XOAI21X1_28 OAI21X1_4/B NAND3X1_3/Y NAND2X1_31/Y gnd OAI21X1_28/Y vdd OAI21X1
XOAI21X1_17 OAI21X1_9/A NAND3X1_2/Y OAI21X1_17/C gnd OAI21X1_17/Y vdd OAI21X1
XFILL_12_1 gnd vdd FILL
XDFFPOSX1_112 NAND2X1_35/A CLKBUF1_4/Y OAI21X1_32/Y gnd vdd DFFPOSX1
XFILL_0_2_1 gnd vdd FILL
XDFFPOSX1_123 NOR2X1_43/A CLKBUF1_5/Y OAI21X1_11/Y gnd vdd DFFPOSX1
XDFFPOSX1_101 INVX1_36/A CLKBUF1_5/Y MUX2X1_26/Y gnd vdd DFFPOSX1
XFILL_16_2_1 gnd vdd FILL
XXNOR2X1_4 XNOR2X1_4/A DFFSR_7/Q gnd DFFSR_7/D vdd XNOR2X1
XINVX1_4 INVX1_4/A gnd INVX1_4/Y vdd INVX1
XFILL_5_1_1 gnd vdd FILL
XFILL_13_0_1 gnd vdd FILL
XDFFSR_8 INVX1_3/A CLKBUF1_3/Y DFFSR_4/R vdd DFFSR_8/D gnd vdd DFFSR
XMUX2X1_27 OAI21X1_6/B INVX1_42/Y NOR2X1_77/Y gnd MUX2X1_27/Y vdd MUX2X1
XMUX2X1_16 INVX4_2/Y INVX1_20/Y MUX2X1_19/S gnd MUX2X1_16/Y vdd MUX2X1
XNAND2X1_42 NAND2X1_42/A NAND3X1_4/Y gnd OAI21X1_39/C vdd NAND2X1
XNAND2X1_53 NAND3X1_5/B NAND3X1_5/C gnd NOR2X1_36/B vdd NAND2X1
XNAND2X1_64 INVX1_9/Y NAND3X1_5/B gnd NAND2X1_64/Y vdd NAND2X1
XNAND2X1_31 NAND2X1_31/A NAND3X1_3/Y gnd NAND2X1_31/Y vdd NAND2X1
XNAND2X1_97 DFFPOSX1_8/Q NAND3X1_15/Y gnd NAND2X1_97/Y vdd NAND2X1
XNAND2X1_75 d_in[1] BUFX4_10/Y gnd OAI21X1_2/B vdd NAND2X1
XNAND2X1_20 AOI21X1_33/A NAND3X1_2/Y gnd OAI21X1_17/C vdd NAND2X1
XNAND2X1_86 AOI21X1_73/B NAND3X1_14/Y gnd NAND2X1_86/Y vdd NAND2X1
XOAI22X1_2 OAI22X1_2/A OAI22X1_2/B OAI22X1_2/C BUFX4_36/Y gnd DFFSR_10/D vdd OAI22X1
XOAI21X1_18 OAI21X1_2/B NAND3X1_2/Y OAI21X1_18/C gnd OAI21X1_18/Y vdd OAI21X1
XOAI21X1_29 MUX2X1_26/A NAND3X1_3/Y OAI21X1_29/C gnd OAI21X1_29/Y vdd OAI21X1
XDFFPOSX1_102 INVX1_42/A CLKBUF1_8/Y MUX2X1_27/Y gnd vdd DFFPOSX1
XDFFPOSX1_124 INVX1_32/A CLKBUF1_4/Y OAI21X1_12/Y gnd vdd DFFPOSX1
XDFFPOSX1_113 AOI21X1_33/A CLKBUF1_11/Y OAI21X1_17/Y gnd vdd DFFPOSX1
XBUFX4_40 DFFSR_1/Q gnd INVX8_2/A vdd BUFX4
XXNOR2X1_5 XNOR2X1_5/A DFFSR_17/Q gnd XNOR2X1_6/A vdd XNOR2X1
XINVX1_5 INVX1_5/A gnd INVX1_5/Y vdd INVX1
.ends

