VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO fifo
  CLASS BLOCK ;
  FOREIGN fifo ;
  ORIGIN 2.600 3.200 ;
  SIZE 210.800 BY 186.400 ;
  PIN vdd
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.200 180.200 205.400 180.800 ;
        RECT 1.400 176.500 1.800 180.200 ;
        RECT 3.800 176.500 4.200 180.200 ;
        RECT 5.400 175.900 5.800 180.200 ;
        RECT 7.000 175.900 7.400 180.200 ;
        RECT 8.600 175.900 9.000 180.200 ;
        RECT 10.200 175.900 10.600 180.200 ;
        RECT 11.800 175.900 12.200 180.200 ;
        RECT 13.400 176.500 13.800 180.200 ;
        RECT 15.800 176.500 16.200 180.200 ;
        RECT 18.200 176.500 18.600 180.200 ;
        RECT 19.800 177.900 20.200 180.200 ;
        RECT 21.400 177.900 21.800 180.200 ;
        RECT 23.000 177.900 23.400 180.200 ;
        RECT 24.600 177.900 25.000 180.200 ;
        RECT 28.600 177.900 29.000 180.200 ;
        RECT 30.200 177.900 30.600 180.200 ;
        RECT 33.400 177.900 33.800 180.200 ;
        RECT 35.000 177.900 35.400 180.200 ;
        RECT 36.600 177.900 37.000 180.200 ;
        RECT 33.300 175.900 33.700 176.000 ;
        RECT 35.000 175.900 35.400 176.200 ;
        RECT 37.400 175.900 37.800 180.200 ;
        RECT 39.000 176.500 39.400 180.200 ;
        RECT 41.400 176.500 41.800 180.200 ;
        RECT 44.600 177.900 45.000 180.200 ;
        RECT 46.200 177.900 46.600 180.200 ;
        RECT 47.800 177.900 48.200 180.200 ;
        RECT 49.400 177.900 49.800 180.200 ;
        RECT 53.400 177.900 53.800 180.200 ;
        RECT 55.000 177.900 55.400 180.200 ;
        RECT 58.200 177.900 58.600 180.200 ;
        RECT 59.800 177.900 60.200 180.200 ;
        RECT 61.400 177.900 61.800 180.200 ;
        RECT 58.100 175.900 58.500 176.000 ;
        RECT 59.800 175.900 60.200 176.200 ;
        RECT 63.000 175.900 63.400 180.200 ;
        RECT 65.800 177.900 66.200 180.200 ;
        RECT 67.400 177.900 67.800 180.200 ;
        RECT 70.200 176.000 70.600 180.200 ;
        RECT 72.600 175.900 73.000 180.200 ;
        RECT 75.400 177.900 75.800 180.200 ;
        RECT 77.000 177.900 77.400 180.200 ;
        RECT 79.800 176.000 80.200 180.200 ;
        RECT 81.400 175.900 81.800 180.200 ;
        RECT 83.000 175.900 83.400 180.200 ;
        RECT 84.600 175.900 85.000 180.200 ;
        RECT 85.400 175.900 85.800 180.200 ;
        RECT 87.000 175.900 87.400 180.200 ;
        RECT 88.600 175.900 89.000 180.200 ;
        RECT 90.200 175.900 90.600 180.200 ;
        RECT 91.800 175.900 92.200 180.200 ;
        RECT 92.600 177.900 93.000 180.200 ;
        RECT 94.200 177.900 94.600 180.200 ;
        RECT 95.800 177.900 96.200 180.200 ;
        RECT 99.000 177.900 99.400 180.200 ;
        RECT 100.600 177.900 101.000 180.200 ;
        RECT 104.600 177.900 105.000 180.200 ;
        RECT 106.200 177.900 106.600 180.200 ;
        RECT 107.800 177.900 108.200 180.200 ;
        RECT 109.400 177.900 109.800 180.200 ;
        RECT 112.600 176.500 113.000 180.200 ;
        RECT 94.200 175.900 94.600 176.200 ;
        RECT 95.800 175.900 96.300 176.000 ;
        RECT 114.200 175.900 114.600 180.200 ;
        RECT 115.000 175.900 115.400 180.200 ;
        RECT 116.600 175.900 117.000 180.200 ;
        RECT 118.200 175.900 118.600 180.200 ;
        RECT 119.800 175.900 120.200 180.200 ;
        RECT 121.400 175.900 121.800 180.200 ;
        RECT 122.200 175.900 122.600 180.200 ;
        RECT 125.400 177.900 125.800 180.200 ;
        RECT 127.800 175.900 128.200 180.200 ;
        RECT 129.400 175.900 129.800 180.200 ;
        RECT 130.200 177.900 130.600 180.200 ;
        RECT 131.800 177.900 132.200 180.200 ;
        RECT 133.400 177.900 133.800 180.200 ;
        RECT 135.000 177.900 135.400 180.200 ;
        RECT 139.000 177.900 139.400 180.200 ;
        RECT 140.600 177.900 141.000 180.200 ;
        RECT 143.800 177.900 144.200 180.200 ;
        RECT 145.400 177.900 145.800 180.200 ;
        RECT 147.000 177.900 147.400 180.200 ;
        RECT 149.400 177.900 149.800 180.200 ;
        RECT 151.000 177.900 151.400 180.200 ;
        RECT 152.600 177.900 153.000 180.200 ;
        RECT 155.800 177.900 156.200 180.200 ;
        RECT 157.400 177.900 157.800 180.200 ;
        RECT 161.400 177.900 161.800 180.200 ;
        RECT 163.000 177.900 163.400 180.200 ;
        RECT 164.600 177.900 165.000 180.200 ;
        RECT 166.200 177.900 166.600 180.200 ;
        RECT 143.700 175.900 144.100 176.000 ;
        RECT 145.400 175.900 145.800 176.200 ;
        RECT 21.900 175.600 35.400 175.900 ;
        RECT 46.700 175.600 60.200 175.900 ;
        RECT 94.200 175.600 107.700 175.900 ;
        RECT 21.900 175.500 22.300 175.600 ;
        RECT 46.700 175.500 47.100 175.600 ;
        RECT 107.300 175.500 107.700 175.600 ;
        RECT 132.300 175.600 145.800 175.900 ;
        RECT 151.000 175.900 151.400 176.200 ;
        RECT 152.700 175.900 153.100 176.000 ;
        RECT 167.000 175.900 167.400 180.200 ;
        RECT 168.600 175.900 169.000 180.200 ;
        RECT 170.200 175.900 170.600 180.200 ;
        RECT 171.800 175.900 172.200 180.200 ;
        RECT 173.400 175.900 173.800 180.200 ;
        RECT 174.200 177.900 174.600 180.200 ;
        RECT 175.800 177.900 176.200 180.200 ;
        RECT 177.400 177.900 177.800 180.200 ;
        RECT 180.600 177.900 181.000 180.200 ;
        RECT 182.200 177.900 182.600 180.200 ;
        RECT 186.200 177.900 186.600 180.200 ;
        RECT 187.800 177.900 188.200 180.200 ;
        RECT 189.400 177.900 189.800 180.200 ;
        RECT 191.000 177.900 191.400 180.200 ;
        RECT 192.600 177.900 193.000 180.200 ;
        RECT 193.400 177.900 193.800 180.200 ;
        RECT 195.000 178.100 195.400 180.200 ;
        RECT 196.600 177.900 197.000 180.200 ;
        RECT 199.000 176.500 199.400 180.200 ;
        RECT 200.600 177.900 201.000 180.200 ;
        RECT 203.000 176.500 203.400 180.200 ;
        RECT 175.800 175.900 176.200 176.200 ;
        RECT 177.500 175.900 177.900 176.000 ;
        RECT 151.000 175.600 164.500 175.900 ;
        RECT 175.800 175.600 189.300 175.900 ;
        RECT 132.300 175.500 132.700 175.600 ;
        RECT 164.100 175.500 164.500 175.600 ;
        RECT 188.900 175.500 189.300 175.600 ;
        RECT 2.700 165.400 3.100 165.500 ;
        RECT 20.300 165.400 20.700 165.500 ;
        RECT 37.900 165.400 38.300 165.500 ;
        RECT 137.100 165.400 137.500 165.500 ;
        RECT 180.100 165.400 180.500 165.500 ;
        RECT 2.700 165.100 16.200 165.400 ;
        RECT 20.300 165.100 33.800 165.400 ;
        RECT 37.900 165.100 51.400 165.400 ;
        RECT 137.100 165.100 150.600 165.400 ;
        RECT 14.100 165.000 14.500 165.100 ;
        RECT 15.800 164.800 16.200 165.100 ;
        RECT 31.700 165.000 32.200 165.100 ;
        RECT 33.400 164.800 33.800 165.100 ;
        RECT 49.300 165.000 49.800 165.100 ;
        RECT 51.000 164.800 51.400 165.100 ;
        RECT 0.600 160.800 1.000 163.100 ;
        RECT 2.200 160.800 2.600 163.100 ;
        RECT 3.800 160.800 4.200 163.100 ;
        RECT 5.400 160.800 5.800 163.100 ;
        RECT 9.400 160.800 9.800 163.100 ;
        RECT 11.000 160.800 11.400 163.100 ;
        RECT 14.200 160.800 14.600 163.100 ;
        RECT 15.800 160.800 16.200 163.100 ;
        RECT 17.400 160.800 17.800 163.100 ;
        RECT 18.200 160.800 18.600 163.100 ;
        RECT 19.800 160.800 20.200 163.100 ;
        RECT 21.400 160.800 21.800 163.100 ;
        RECT 23.000 160.800 23.400 163.100 ;
        RECT 27.000 160.800 27.400 163.100 ;
        RECT 28.600 160.800 29.000 163.100 ;
        RECT 31.800 160.800 32.200 163.100 ;
        RECT 33.400 160.800 33.800 163.100 ;
        RECT 35.000 160.800 35.400 163.100 ;
        RECT 35.800 160.800 36.200 163.100 ;
        RECT 37.400 160.800 37.800 163.100 ;
        RECT 39.000 160.800 39.400 163.100 ;
        RECT 40.600 160.800 41.000 163.100 ;
        RECT 44.600 160.800 45.000 163.100 ;
        RECT 46.200 160.800 46.600 163.100 ;
        RECT 49.400 160.800 49.800 163.100 ;
        RECT 51.000 160.800 51.400 163.100 ;
        RECT 52.600 160.800 53.000 163.100 ;
        RECT 55.000 160.800 55.400 165.100 ;
        RECT 56.600 160.800 57.000 164.500 ;
        RECT 58.200 160.800 58.600 165.100 ;
        RECT 60.300 160.800 60.700 163.100 ;
        RECT 61.400 160.800 61.800 163.100 ;
        RECT 63.000 160.800 63.400 163.100 ;
        RECT 64.600 160.800 65.000 164.500 ;
        RECT 68.600 160.800 69.000 165.100 ;
        RECT 70.200 160.800 70.600 165.000 ;
        RECT 73.000 160.800 73.400 163.100 ;
        RECT 74.600 160.800 75.000 163.100 ;
        RECT 77.400 160.800 77.800 165.100 ;
        RECT 79.000 160.800 79.400 165.100 ;
        RECT 81.100 160.800 81.500 163.100 ;
        RECT 82.200 160.800 82.600 163.100 ;
        RECT 83.800 160.800 84.200 163.100 ;
        RECT 85.400 160.800 85.800 165.100 ;
        RECT 88.200 160.800 88.600 163.100 ;
        RECT 89.800 160.800 90.200 163.100 ;
        RECT 92.600 160.800 93.000 165.000 ;
        RECT 95.000 161.100 95.500 164.400 ;
        RECT 95.100 160.800 95.500 161.100 ;
        RECT 98.100 160.800 98.600 164.400 ;
        RECT 100.600 160.800 101.000 165.100 ;
        RECT 104.600 160.800 105.000 165.100 ;
        RECT 105.400 160.800 105.800 163.100 ;
        RECT 107.000 160.800 107.400 163.100 ;
        RECT 109.400 160.800 109.800 165.100 ;
        RECT 111.800 160.800 112.200 165.100 ;
        RECT 112.600 160.800 113.000 163.100 ;
        RECT 114.200 160.800 114.600 163.100 ;
        RECT 115.000 160.800 115.400 163.100 ;
        RECT 116.600 160.800 117.000 162.900 ;
        RECT 118.200 160.800 118.600 165.100 ;
        RECT 120.300 160.800 120.700 163.100 ;
        RECT 121.400 160.800 121.800 165.100 ;
        RECT 123.800 160.800 124.200 165.100 ;
        RECT 126.500 160.800 126.900 163.100 ;
        RECT 128.600 160.800 129.000 165.100 ;
        RECT 148.500 165.000 148.900 165.100 ;
        RECT 150.200 164.800 150.600 165.100 ;
        RECT 167.000 165.100 180.500 165.400 ;
        RECT 167.000 164.800 167.400 165.100 ;
        RECT 168.700 165.000 169.100 165.100 ;
        RECT 130.200 161.100 130.700 164.400 ;
        RECT 130.300 160.800 130.700 161.100 ;
        RECT 133.300 160.800 133.800 164.400 ;
        RECT 135.000 160.800 135.400 163.100 ;
        RECT 136.600 160.800 137.000 163.100 ;
        RECT 138.200 160.800 138.600 163.100 ;
        RECT 139.800 160.800 140.200 163.100 ;
        RECT 143.800 160.800 144.200 163.100 ;
        RECT 145.400 160.800 145.800 163.100 ;
        RECT 148.600 160.800 149.000 163.100 ;
        RECT 150.200 160.800 150.600 163.100 ;
        RECT 151.800 160.800 152.200 163.100 ;
        RECT 155.000 160.800 155.500 164.400 ;
        RECT 158.100 161.100 158.600 164.400 ;
        RECT 160.600 161.100 161.100 164.400 ;
        RECT 158.100 160.800 158.500 161.100 ;
        RECT 160.700 160.800 161.100 161.100 ;
        RECT 163.700 160.800 164.200 164.400 ;
        RECT 165.400 160.800 165.800 163.100 ;
        RECT 167.000 160.800 167.400 163.100 ;
        RECT 168.600 160.800 169.000 163.100 ;
        RECT 171.800 160.800 172.200 163.100 ;
        RECT 173.400 160.800 173.800 163.100 ;
        RECT 177.400 160.800 177.800 163.100 ;
        RECT 179.000 160.800 179.400 163.100 ;
        RECT 180.600 160.800 181.000 163.100 ;
        RECT 182.200 160.800 182.600 163.100 ;
        RECT 183.000 160.800 183.400 163.100 ;
        RECT 184.600 160.800 185.000 163.100 ;
        RECT 185.700 160.800 186.100 163.100 ;
        RECT 187.800 160.800 188.200 165.100 ;
        RECT 189.400 160.800 189.800 164.500 ;
        RECT 192.600 161.100 193.100 164.400 ;
        RECT 192.700 160.800 193.100 161.100 ;
        RECT 195.700 160.800 196.200 164.400 ;
        RECT 197.400 160.800 197.800 165.100 ;
        RECT 199.500 160.800 199.900 163.100 ;
        RECT 200.600 160.800 201.000 163.100 ;
        RECT 202.200 160.800 202.600 162.900 ;
        RECT 204.600 160.800 205.000 163.100 ;
        RECT 0.200 160.200 205.400 160.800 ;
        RECT 1.400 156.500 1.800 160.200 ;
        RECT 3.800 156.500 4.200 160.200 ;
        RECT 6.200 156.000 6.600 160.200 ;
        RECT 9.000 157.900 9.400 160.200 ;
        RECT 10.600 157.900 11.000 160.200 ;
        RECT 13.400 155.900 13.800 160.200 ;
        RECT 15.000 155.900 15.400 160.200 ;
        RECT 17.400 157.900 17.800 160.200 ;
        RECT 19.000 157.900 19.400 160.200 ;
        RECT 20.600 157.900 21.000 160.200 ;
        RECT 22.200 157.900 22.600 160.200 ;
        RECT 26.200 157.900 26.600 160.200 ;
        RECT 27.800 157.900 28.200 160.200 ;
        RECT 31.000 157.900 31.400 160.200 ;
        RECT 32.600 157.900 33.000 160.200 ;
        RECT 34.200 157.900 34.600 160.200 ;
        RECT 35.800 156.500 36.200 160.200 ;
        RECT 30.900 155.900 31.300 156.000 ;
        RECT 32.600 155.900 33.000 156.200 ;
        RECT 39.800 155.900 40.200 160.200 ;
        RECT 41.400 156.000 41.800 160.200 ;
        RECT 44.200 157.900 44.600 160.200 ;
        RECT 45.800 157.900 46.200 160.200 ;
        RECT 48.600 155.900 49.000 160.200 ;
        RECT 51.800 155.900 52.200 160.200 ;
        RECT 53.900 157.900 54.300 160.200 ;
        RECT 55.000 157.900 55.400 160.200 ;
        RECT 56.600 157.900 57.000 160.200 ;
        RECT 58.200 156.500 58.600 160.200 ;
        RECT 61.400 156.000 61.800 160.200 ;
        RECT 64.200 157.900 64.600 160.200 ;
        RECT 65.800 157.900 66.200 160.200 ;
        RECT 68.600 155.900 69.000 160.200 ;
        RECT 70.200 155.900 70.600 160.200 ;
        RECT 72.300 157.900 72.700 160.200 ;
        RECT 73.400 157.900 73.800 160.200 ;
        RECT 75.000 157.900 75.400 160.200 ;
        RECT 75.800 157.900 76.200 160.200 ;
        RECT 77.400 157.900 77.800 160.200 ;
        RECT 78.200 157.900 78.600 160.200 ;
        RECT 79.800 157.900 80.200 160.200 ;
        RECT 81.400 157.900 81.800 160.200 ;
        RECT 84.600 157.900 85.000 160.200 ;
        RECT 86.200 157.900 86.600 160.200 ;
        RECT 90.200 157.900 90.600 160.200 ;
        RECT 91.800 157.900 92.200 160.200 ;
        RECT 93.400 157.900 93.800 160.200 ;
        RECT 95.000 157.900 95.400 160.200 ;
        RECT 96.100 157.900 96.500 160.200 ;
        RECT 79.800 155.900 80.200 156.200 ;
        RECT 81.500 155.900 81.900 156.000 ;
        RECT 98.200 155.900 98.600 160.200 ;
        RECT 100.600 155.900 101.000 160.200 ;
        RECT 103.000 157.900 103.400 160.200 ;
        RECT 104.600 155.900 105.000 160.200 ;
        RECT 107.000 157.900 107.400 160.200 ;
        RECT 108.600 157.900 109.000 160.200 ;
        RECT 109.400 155.900 109.800 160.200 ;
        RECT 112.600 156.500 113.000 160.200 ;
        RECT 114.200 155.900 114.600 160.200 ;
        RECT 115.000 157.900 115.400 160.200 ;
        RECT 116.600 157.900 117.000 160.200 ;
        RECT 117.400 155.900 117.800 160.200 ;
        RECT 119.800 157.900 120.200 160.200 ;
        RECT 121.400 157.900 121.800 160.200 ;
        RECT 122.200 157.900 122.600 160.200 ;
        RECT 123.800 157.900 124.200 160.200 ;
        RECT 124.600 157.900 125.000 160.200 ;
        RECT 126.200 157.900 126.600 160.200 ;
        RECT 127.800 157.900 128.200 160.200 ;
        RECT 129.400 157.900 129.800 160.200 ;
        RECT 133.400 157.900 133.800 160.200 ;
        RECT 135.000 157.900 135.400 160.200 ;
        RECT 138.200 157.900 138.600 160.200 ;
        RECT 139.800 157.900 140.200 160.200 ;
        RECT 141.400 157.900 141.800 160.200 ;
        RECT 142.200 157.900 142.600 160.200 ;
        RECT 143.800 157.900 144.200 160.200 ;
        RECT 145.400 157.900 145.800 160.200 ;
        RECT 147.000 157.900 147.400 160.200 ;
        RECT 151.000 157.900 151.400 160.200 ;
        RECT 152.600 157.900 153.000 160.200 ;
        RECT 155.800 157.900 156.200 160.200 ;
        RECT 157.400 157.900 157.800 160.200 ;
        RECT 159.000 157.900 159.400 160.200 ;
        RECT 161.400 157.900 161.800 160.200 ;
        RECT 163.000 157.900 163.400 160.200 ;
        RECT 164.600 157.900 165.000 160.200 ;
        RECT 167.800 157.900 168.200 160.200 ;
        RECT 169.400 157.900 169.800 160.200 ;
        RECT 173.400 157.900 173.800 160.200 ;
        RECT 175.000 157.900 175.400 160.200 ;
        RECT 176.600 157.900 177.000 160.200 ;
        RECT 178.200 157.900 178.600 160.200 ;
        RECT 138.100 155.900 138.500 156.000 ;
        RECT 139.800 155.900 140.200 156.200 ;
        RECT 155.700 155.900 156.100 156.000 ;
        RECT 157.400 155.900 157.800 156.200 ;
        RECT 19.500 155.600 33.000 155.900 ;
        RECT 79.800 155.600 93.300 155.900 ;
        RECT 19.500 155.500 19.900 155.600 ;
        RECT 92.900 155.500 93.300 155.600 ;
        RECT 126.700 155.600 140.200 155.900 ;
        RECT 144.300 155.600 157.800 155.900 ;
        RECT 163.000 155.900 163.400 156.200 ;
        RECT 164.700 155.900 165.100 156.000 ;
        RECT 180.600 155.900 181.000 160.200 ;
        RECT 183.000 155.900 183.400 160.200 ;
        RECT 183.800 155.900 184.200 160.200 ;
        RECT 185.900 157.900 186.300 160.200 ;
        RECT 187.000 157.900 187.400 160.200 ;
        RECT 188.600 155.900 189.000 160.200 ;
        RECT 190.700 157.900 191.100 160.200 ;
        RECT 192.600 156.100 193.000 160.200 ;
        RECT 194.200 157.900 194.600 160.200 ;
        RECT 195.800 156.000 196.200 160.200 ;
        RECT 198.600 157.900 199.000 160.200 ;
        RECT 200.200 157.900 200.600 160.200 ;
        RECT 203.000 155.900 203.400 160.200 ;
        RECT 163.000 155.600 176.500 155.900 ;
        RECT 126.700 155.500 127.100 155.600 ;
        RECT 144.300 155.500 144.700 155.600 ;
        RECT 176.100 155.500 176.500 155.600 ;
        RECT 69.100 145.400 69.500 145.500 ;
        RECT 69.100 145.100 82.600 145.400 ;
        RECT 1.400 140.800 1.800 145.000 ;
        RECT 4.200 140.800 4.600 143.100 ;
        RECT 5.800 140.800 6.200 143.100 ;
        RECT 8.600 140.800 9.000 145.100 ;
        RECT 10.200 140.800 10.600 145.100 ;
        RECT 12.300 140.800 12.700 143.100 ;
        RECT 14.200 140.800 14.600 144.500 ;
        RECT 16.600 140.800 17.000 143.100 ;
        RECT 18.200 140.800 18.600 143.100 ;
        RECT 19.300 140.800 19.700 143.100 ;
        RECT 21.400 140.800 21.800 145.100 ;
        RECT 23.000 140.800 23.400 145.000 ;
        RECT 25.800 140.800 26.200 143.100 ;
        RECT 27.400 140.800 27.800 143.100 ;
        RECT 30.200 140.800 30.600 145.100 ;
        RECT 32.600 140.800 33.000 145.000 ;
        RECT 35.400 140.800 35.800 143.100 ;
        RECT 37.000 140.800 37.400 143.100 ;
        RECT 39.800 140.800 40.200 145.100 ;
        RECT 42.200 140.800 42.600 145.000 ;
        RECT 45.000 140.800 45.400 143.100 ;
        RECT 46.600 140.800 47.000 143.100 ;
        RECT 49.400 140.800 49.800 145.100 ;
        RECT 53.400 140.800 53.800 143.100 ;
        RECT 54.200 140.800 54.600 143.100 ;
        RECT 55.800 140.800 56.200 143.100 ;
        RECT 56.900 140.800 57.300 143.100 ;
        RECT 59.000 140.800 59.400 145.100 ;
        RECT 60.600 140.800 61.000 144.500 ;
        RECT 62.200 140.800 62.600 145.100 ;
        RECT 63.000 140.800 63.400 143.100 ;
        RECT 66.200 140.800 66.600 145.100 ;
        RECT 80.500 145.000 81.000 145.100 ;
        RECT 82.200 144.800 82.600 145.100 ;
        RECT 67.000 140.800 67.400 143.100 ;
        RECT 68.600 140.800 69.000 143.100 ;
        RECT 70.200 140.800 70.600 143.100 ;
        RECT 71.800 140.800 72.200 143.100 ;
        RECT 75.800 140.800 76.200 143.100 ;
        RECT 77.400 140.800 77.800 143.100 ;
        RECT 80.600 140.800 81.000 143.100 ;
        RECT 82.200 140.800 82.600 143.100 ;
        RECT 83.800 140.800 84.200 143.100 ;
        RECT 84.600 140.800 85.000 143.100 ;
        RECT 86.200 140.800 86.600 145.100 ;
        RECT 88.300 140.800 88.700 143.100 ;
        RECT 89.400 140.800 89.800 143.100 ;
        RECT 91.000 140.800 91.400 143.100 ;
        RECT 92.600 140.800 93.000 145.100 ;
        RECT 95.400 140.800 95.800 143.100 ;
        RECT 97.000 140.800 97.400 143.100 ;
        RECT 99.800 140.800 100.200 145.000 ;
        RECT 103.800 140.800 104.200 142.900 ;
        RECT 105.400 140.800 105.800 143.100 ;
        RECT 106.200 140.800 106.600 143.100 ;
        RECT 107.800 140.800 108.200 142.900 ;
        RECT 111.000 140.800 111.400 145.100 ;
        RECT 111.800 140.800 112.200 143.100 ;
        RECT 113.400 140.800 113.800 143.100 ;
        RECT 114.200 140.800 114.600 143.100 ;
        RECT 115.800 140.800 116.200 142.900 ;
        RECT 117.400 140.800 117.800 143.100 ;
        RECT 119.000 140.800 119.400 142.900 ;
        RECT 120.600 140.800 121.000 143.100 ;
        RECT 122.200 140.800 122.600 142.900 ;
        RECT 123.800 140.800 124.200 143.100 ;
        RECT 125.400 140.800 125.800 142.900 ;
        RECT 127.000 140.800 127.400 143.100 ;
        RECT 128.600 140.800 129.000 142.900 ;
        RECT 130.200 140.800 130.600 145.100 ;
        RECT 132.600 140.800 133.000 145.100 ;
        RECT 134.200 140.800 134.600 144.500 ;
        RECT 135.800 140.800 136.200 145.100 ;
        RECT 139.000 140.800 139.500 144.400 ;
        RECT 142.100 141.100 142.600 144.400 ;
        RECT 142.100 140.800 142.500 141.100 ;
        RECT 143.800 140.800 144.200 143.100 ;
        RECT 145.400 140.800 145.800 143.100 ;
        RECT 146.200 140.800 146.600 143.100 ;
        RECT 147.800 140.800 148.200 143.100 ;
        RECT 149.400 140.800 149.800 144.500 ;
        RECT 155.800 140.800 156.200 144.500 ;
        RECT 157.700 140.800 158.100 143.100 ;
        RECT 159.800 140.800 160.200 145.100 ;
        RECT 160.600 140.800 161.000 143.100 ;
        RECT 162.200 140.800 162.600 143.100 ;
        RECT 163.800 140.800 164.200 143.100 ;
        RECT 164.600 140.800 165.000 145.100 ;
        RECT 166.700 140.800 167.100 143.100 ;
        RECT 170.200 140.800 170.600 144.500 ;
        RECT 171.800 140.800 172.200 143.100 ;
        RECT 173.400 140.800 173.800 143.100 ;
        RECT 175.800 140.800 176.200 144.500 ;
        RECT 177.400 140.800 177.800 143.100 ;
        RECT 179.000 140.800 179.400 143.100 ;
        RECT 181.400 140.800 181.800 145.100 ;
        RECT 183.000 140.800 183.400 144.500 ;
        RECT 187.800 140.800 188.200 145.100 ;
        RECT 188.600 140.800 189.000 143.100 ;
        RECT 190.200 140.800 190.600 143.100 ;
        RECT 191.000 140.800 191.400 145.100 ;
        RECT 193.400 140.800 193.800 143.100 ;
        RECT 195.000 140.800 195.400 142.900 ;
        RECT 197.400 140.800 197.800 142.900 ;
        RECT 199.000 140.800 199.400 143.100 ;
        RECT 200.600 140.800 201.000 144.900 ;
        RECT 202.200 140.800 202.600 143.100 ;
        RECT 203.800 140.800 204.200 144.500 ;
        RECT 0.200 140.200 205.400 140.800 ;
        RECT 0.600 137.900 1.000 140.200 ;
        RECT 2.200 137.900 2.600 140.200 ;
        RECT 3.800 137.900 4.200 140.200 ;
        RECT 5.400 137.900 5.800 140.200 ;
        RECT 9.400 137.900 9.800 140.200 ;
        RECT 11.000 137.900 11.400 140.200 ;
        RECT 14.200 137.900 14.600 140.200 ;
        RECT 15.800 137.900 16.200 140.200 ;
        RECT 17.400 137.900 17.800 140.200 ;
        RECT 18.200 137.900 18.600 140.200 ;
        RECT 19.800 137.900 20.200 140.200 ;
        RECT 20.600 137.900 21.000 140.200 ;
        RECT 22.200 137.900 22.600 140.200 ;
        RECT 23.800 137.900 24.200 140.200 ;
        RECT 25.400 137.900 25.800 140.200 ;
        RECT 29.400 137.900 29.800 140.200 ;
        RECT 31.000 137.900 31.400 140.200 ;
        RECT 34.200 137.900 34.600 140.200 ;
        RECT 35.800 137.900 36.200 140.200 ;
        RECT 37.400 137.900 37.800 140.200 ;
        RECT 14.100 135.900 14.500 136.000 ;
        RECT 15.800 135.900 16.200 136.200 ;
        RECT 34.100 135.900 34.500 136.000 ;
        RECT 35.800 135.900 36.200 136.200 ;
        RECT 38.200 135.900 38.600 140.200 ;
        RECT 40.300 137.900 40.700 140.200 ;
        RECT 42.200 136.500 42.600 140.200 ;
        RECT 44.900 137.900 45.300 140.200 ;
        RECT 47.000 135.900 47.400 140.200 ;
        RECT 49.400 136.500 49.800 140.200 ;
        RECT 53.400 136.000 53.800 140.200 ;
        RECT 56.200 137.900 56.600 140.200 ;
        RECT 57.800 137.900 58.200 140.200 ;
        RECT 60.600 135.900 61.000 140.200 ;
        RECT 62.200 137.900 62.600 140.200 ;
        RECT 63.800 137.900 64.200 140.200 ;
        RECT 64.900 137.900 65.300 140.200 ;
        RECT 67.000 135.900 67.400 140.200 ;
        RECT 67.800 135.900 68.200 140.200 ;
        RECT 69.900 137.900 70.300 140.200 ;
        RECT 71.000 137.900 71.400 140.200 ;
        RECT 72.600 137.900 73.000 140.200 ;
        RECT 74.200 136.500 74.600 140.200 ;
        RECT 76.600 137.900 77.000 140.200 ;
        RECT 78.200 137.900 78.600 140.200 ;
        RECT 79.300 137.900 79.700 140.200 ;
        RECT 81.400 135.900 81.800 140.200 ;
        RECT 83.000 135.900 83.400 140.200 ;
        RECT 85.800 137.900 86.200 140.200 ;
        RECT 87.400 137.900 87.800 140.200 ;
        RECT 90.200 136.000 90.600 140.200 ;
        RECT 91.800 137.900 92.200 140.200 ;
        RECT 93.400 137.900 93.800 140.200 ;
        RECT 94.500 137.900 94.900 140.200 ;
        RECT 96.600 135.900 97.000 140.200 ;
        RECT 97.400 135.900 97.800 140.200 ;
        RECT 99.000 136.500 99.400 140.200 ;
        RECT 103.000 136.500 103.400 140.200 ;
        RECT 104.600 135.900 105.000 140.200 ;
        RECT 106.200 136.100 106.600 140.200 ;
        RECT 108.800 135.900 109.200 140.200 ;
        RECT 110.200 135.900 110.600 140.200 ;
        RECT 112.300 137.900 112.700 140.200 ;
        RECT 113.400 137.900 113.800 140.200 ;
        RECT 115.000 137.900 115.400 140.200 ;
        RECT 116.600 135.900 117.000 140.200 ;
        RECT 119.400 137.900 119.800 140.200 ;
        RECT 121.000 137.900 121.400 140.200 ;
        RECT 123.800 136.000 124.200 140.200 ;
        RECT 125.400 137.900 125.800 140.200 ;
        RECT 127.000 137.900 127.400 140.200 ;
        RECT 127.800 137.900 128.200 140.200 ;
        RECT 129.400 137.900 129.800 140.200 ;
        RECT 130.200 135.900 130.600 140.200 ;
        RECT 132.600 135.900 133.000 140.200 ;
        RECT 135.000 135.900 135.400 140.200 ;
        RECT 139.000 136.500 139.400 140.200 ;
        RECT 140.600 135.900 141.000 140.200 ;
        RECT 142.200 136.500 142.600 140.200 ;
        RECT 144.600 136.500 145.000 140.200 ;
        RECT 146.200 135.900 146.600 140.200 ;
        RECT 147.800 136.500 148.200 140.200 ;
        RECT 149.400 135.900 149.800 140.200 ;
        RECT 152.600 136.000 153.000 140.200 ;
        RECT 155.400 137.900 155.800 140.200 ;
        RECT 157.000 137.900 157.400 140.200 ;
        RECT 159.800 135.900 160.200 140.200 ;
        RECT 163.000 135.900 163.400 140.200 ;
        RECT 163.800 137.900 164.200 140.200 ;
        RECT 166.200 136.100 166.600 140.200 ;
        RECT 168.800 135.900 169.200 140.200 ;
        RECT 170.200 137.900 170.600 140.200 ;
        RECT 171.800 137.900 172.200 140.200 ;
        RECT 172.900 137.900 173.300 140.200 ;
        RECT 175.000 135.900 175.400 140.200 ;
        RECT 176.600 138.100 177.000 140.200 ;
        RECT 178.200 137.900 178.600 140.200 ;
        RECT 179.000 137.900 179.400 140.200 ;
        RECT 180.600 137.900 181.000 140.200 ;
        RECT 182.200 136.100 182.600 140.200 ;
        RECT 183.800 137.900 184.200 140.200 ;
        RECT 184.900 137.900 185.300 140.200 ;
        RECT 187.000 135.900 187.400 140.200 ;
        RECT 187.800 137.900 188.200 140.200 ;
        RECT 189.400 137.900 189.800 140.200 ;
        RECT 190.200 137.900 190.600 140.200 ;
        RECT 191.800 137.900 192.200 140.200 ;
        RECT 193.400 138.100 193.800 140.200 ;
        RECT 195.000 137.900 195.400 140.200 ;
        RECT 197.400 136.500 197.800 140.200 ;
        RECT 199.800 136.600 200.300 140.200 ;
        RECT 202.900 139.900 203.300 140.200 ;
        RECT 202.900 136.600 203.400 139.900 ;
        RECT 2.700 135.600 16.200 135.900 ;
        RECT 22.700 135.600 36.200 135.900 ;
        RECT 2.700 135.500 3.100 135.600 ;
        RECT 22.700 135.500 23.100 135.600 ;
        RECT 1.400 120.800 1.800 125.000 ;
        RECT 4.200 120.800 4.600 123.100 ;
        RECT 5.800 120.800 6.200 123.100 ;
        RECT 8.600 120.800 9.000 125.100 ;
        RECT 10.200 120.800 10.600 123.100 ;
        RECT 12.400 120.800 12.800 125.100 ;
        RECT 15.000 120.800 15.400 124.900 ;
        RECT 17.400 120.800 17.800 125.000 ;
        RECT 20.200 120.800 20.600 123.100 ;
        RECT 21.800 120.800 22.200 123.100 ;
        RECT 24.600 120.800 25.000 125.100 ;
        RECT 26.200 120.800 26.600 125.100 ;
        RECT 28.300 120.800 28.700 123.100 ;
        RECT 29.400 120.800 29.800 123.100 ;
        RECT 31.000 120.800 31.400 123.100 ;
        RECT 32.600 120.800 33.000 125.000 ;
        RECT 35.400 120.800 35.800 123.100 ;
        RECT 37.000 120.800 37.400 123.100 ;
        RECT 39.800 120.800 40.200 125.100 ;
        RECT 41.400 120.800 41.800 123.100 ;
        RECT 43.000 120.800 43.400 123.100 ;
        RECT 43.800 120.800 44.200 125.100 ;
        RECT 45.900 120.800 46.300 123.100 ;
        RECT 47.000 120.800 47.400 125.100 ;
        RECT 50.200 120.800 50.600 125.100 ;
        RECT 53.400 120.800 53.800 124.500 ;
        RECT 56.100 120.800 56.500 123.100 ;
        RECT 58.200 120.800 58.600 125.100 ;
        RECT 59.000 120.800 59.400 123.100 ;
        RECT 60.600 120.800 61.000 123.100 ;
        RECT 61.400 120.800 61.800 123.100 ;
        RECT 63.300 120.800 63.700 123.100 ;
        RECT 65.400 120.800 65.800 125.100 ;
        RECT 66.200 120.800 66.600 125.100 ;
        RECT 68.300 120.800 68.700 123.100 ;
        RECT 69.400 120.800 69.800 125.100 ;
        RECT 71.500 120.800 71.900 123.100 ;
        RECT 73.400 120.800 73.800 125.100 ;
        RECT 76.200 120.800 76.600 123.100 ;
        RECT 77.800 120.800 78.200 123.100 ;
        RECT 80.600 120.800 81.000 125.000 ;
        RECT 82.500 120.800 82.900 123.100 ;
        RECT 84.600 120.800 85.000 125.100 ;
        RECT 87.000 120.800 87.400 125.100 ;
        RECT 88.600 120.800 89.000 123.100 ;
        RECT 90.200 120.800 90.600 125.100 ;
        RECT 93.000 120.800 93.400 123.100 ;
        RECT 94.600 120.800 95.000 123.100 ;
        RECT 97.400 120.800 97.800 125.000 ;
        RECT 99.000 120.800 99.400 123.100 ;
        RECT 100.600 120.800 101.000 123.100 ;
        RECT 103.300 120.800 103.700 123.100 ;
        RECT 105.400 120.800 105.800 125.100 ;
        RECT 106.500 120.800 106.900 123.100 ;
        RECT 108.600 120.800 109.000 125.100 ;
        RECT 109.400 120.800 109.800 125.100 ;
        RECT 112.600 120.800 113.000 125.100 ;
        RECT 115.000 120.800 115.400 125.100 ;
        RECT 115.800 120.800 116.200 125.100 ;
        RECT 119.000 120.800 119.400 125.100 ;
        RECT 121.800 120.800 122.200 123.100 ;
        RECT 123.400 120.800 123.800 123.100 ;
        RECT 126.200 120.800 126.600 125.000 ;
        RECT 128.600 120.800 129.000 125.000 ;
        RECT 131.400 120.800 131.800 123.100 ;
        RECT 133.000 120.800 133.400 123.100 ;
        RECT 135.800 120.800 136.200 125.100 ;
        RECT 137.400 120.800 137.800 125.100 ;
        RECT 139.500 120.800 139.900 123.100 ;
        RECT 140.600 120.800 141.000 123.100 ;
        RECT 142.200 120.800 142.600 123.100 ;
        RECT 143.000 120.800 143.400 123.100 ;
        RECT 145.400 120.800 145.800 125.100 ;
        RECT 148.200 120.800 148.600 123.100 ;
        RECT 149.800 120.800 150.200 123.100 ;
        RECT 152.600 120.800 153.000 125.000 ;
        RECT 155.800 120.800 156.200 125.100 ;
        RECT 159.800 120.800 160.200 124.500 ;
        RECT 163.000 120.800 163.400 124.500 ;
        RECT 164.900 120.800 165.300 123.100 ;
        RECT 167.000 120.800 167.400 125.100 ;
        RECT 168.600 120.800 169.000 124.500 ;
        RECT 171.300 120.800 171.700 123.100 ;
        RECT 173.400 120.800 173.800 125.100 ;
        RECT 175.000 120.800 175.400 124.500 ;
        RECT 176.600 120.800 177.000 125.100 ;
        RECT 177.400 120.800 177.800 123.100 ;
        RECT 179.000 120.800 179.400 123.100 ;
        RECT 179.800 120.800 180.200 123.100 ;
        RECT 181.400 120.800 181.800 123.100 ;
        RECT 183.000 120.800 183.400 124.500 ;
        RECT 184.600 120.800 185.000 125.100 ;
        RECT 185.400 120.800 185.800 125.100 ;
        RECT 187.000 120.800 187.400 125.100 ;
        RECT 187.800 120.800 188.200 125.100 ;
        RECT 189.400 120.800 189.800 125.100 ;
        RECT 190.200 120.800 190.600 125.100 ;
        RECT 191.800 120.800 192.200 125.100 ;
        RECT 193.400 120.800 193.800 124.900 ;
        RECT 196.000 120.800 196.400 125.100 ;
        RECT 198.200 120.800 198.600 124.500 ;
        RECT 201.400 120.800 201.800 123.100 ;
        RECT 202.200 120.800 202.600 125.100 ;
        RECT 0.200 120.200 205.400 120.800 ;
        RECT 1.400 116.000 1.800 120.200 ;
        RECT 4.200 117.900 4.600 120.200 ;
        RECT 5.800 117.900 6.200 120.200 ;
        RECT 8.600 115.900 9.000 120.200 ;
        RECT 11.000 116.000 11.400 120.200 ;
        RECT 13.800 117.900 14.200 120.200 ;
        RECT 15.400 117.900 15.800 120.200 ;
        RECT 18.200 115.900 18.600 120.200 ;
        RECT 19.800 117.900 20.200 120.200 ;
        RECT 22.200 116.100 22.600 120.200 ;
        RECT 24.800 115.900 25.200 120.200 ;
        RECT 27.000 116.000 27.400 120.200 ;
        RECT 29.800 117.900 30.200 120.200 ;
        RECT 31.400 117.900 31.800 120.200 ;
        RECT 34.200 115.900 34.600 120.200 ;
        RECT 35.800 117.900 36.200 120.200 ;
        RECT 37.400 117.900 37.800 120.200 ;
        RECT 38.500 117.900 38.900 120.200 ;
        RECT 40.600 115.900 41.000 120.200 ;
        RECT 41.400 115.900 41.800 120.200 ;
        RECT 43.500 117.900 43.900 120.200 ;
        RECT 46.200 116.500 46.600 120.200 ;
        RECT 47.800 115.900 48.200 120.200 ;
        RECT 49.400 116.500 49.800 120.200 ;
        RECT 52.600 115.900 53.000 120.200 ;
        RECT 54.700 117.900 55.100 120.200 ;
        RECT 55.800 117.900 56.200 120.200 ;
        RECT 57.400 117.900 57.800 120.200 ;
        RECT 59.800 116.500 60.200 120.200 ;
        RECT 61.400 115.900 61.800 120.200 ;
        RECT 63.500 117.900 63.900 120.200 ;
        RECT 65.400 115.900 65.800 120.200 ;
        RECT 68.200 117.900 68.600 120.200 ;
        RECT 69.800 117.900 70.200 120.200 ;
        RECT 72.600 116.000 73.000 120.200 ;
        RECT 74.200 115.900 74.600 120.200 ;
        RECT 75.800 116.500 76.200 120.200 ;
        RECT 78.200 116.500 78.600 120.200 ;
        RECT 79.800 115.900 80.200 120.200 ;
        RECT 81.400 116.500 81.800 120.200 ;
        RECT 83.000 115.900 83.400 120.200 ;
        RECT 85.400 116.500 85.800 120.200 ;
        RECT 87.000 115.900 87.400 120.200 ;
        RECT 89.100 117.900 89.500 120.200 ;
        RECT 90.200 117.900 90.600 120.200 ;
        RECT 91.800 117.900 92.200 120.200 ;
        RECT 93.400 116.000 93.800 120.200 ;
        RECT 96.200 117.900 96.600 120.200 ;
        RECT 97.800 117.900 98.200 120.200 ;
        RECT 100.600 115.900 101.000 120.200 ;
        RECT 103.800 117.900 104.200 120.200 ;
        RECT 105.400 117.900 105.800 120.200 ;
        RECT 106.500 117.900 106.900 120.200 ;
        RECT 108.600 115.900 109.000 120.200 ;
        RECT 110.200 116.500 110.600 120.200 ;
        RECT 111.800 115.900 112.200 120.200 ;
        RECT 113.400 116.600 113.900 120.200 ;
        RECT 116.500 119.900 116.900 120.200 ;
        RECT 116.500 116.600 117.000 119.900 ;
        RECT 118.200 115.900 118.600 120.200 ;
        RECT 119.800 116.500 120.200 120.200 ;
        RECT 121.700 117.900 122.100 120.200 ;
        RECT 123.800 115.900 124.200 120.200 ;
        RECT 125.400 116.500 125.800 120.200 ;
        RECT 128.100 117.900 128.500 120.200 ;
        RECT 130.200 115.900 130.600 120.200 ;
        RECT 131.000 117.900 131.400 120.200 ;
        RECT 132.600 117.900 133.000 120.200 ;
        RECT 133.400 117.900 133.800 120.200 ;
        RECT 135.000 117.900 135.400 120.200 ;
        RECT 136.600 117.900 137.000 120.200 ;
        RECT 138.200 117.900 138.600 120.200 ;
        RECT 142.200 117.900 142.600 120.200 ;
        RECT 143.800 117.900 144.200 120.200 ;
        RECT 147.000 117.900 147.400 120.200 ;
        RECT 148.600 117.900 149.000 120.200 ;
        RECT 150.200 117.900 150.600 120.200 ;
        RECT 146.900 115.900 147.400 116.000 ;
        RECT 148.600 115.900 149.000 116.200 ;
        RECT 152.600 115.900 153.000 120.200 ;
        RECT 156.600 116.500 157.000 120.200 ;
        RECT 159.800 116.500 160.200 120.200 ;
        RECT 162.200 118.100 162.600 120.200 ;
        RECT 163.800 117.900 164.200 120.200 ;
        RECT 164.600 115.900 165.000 120.200 ;
        RECT 166.700 117.900 167.100 120.200 ;
        RECT 167.800 117.900 168.200 120.200 ;
        RECT 169.400 117.900 169.800 120.200 ;
        RECT 171.000 117.900 171.400 120.200 ;
        RECT 174.200 117.900 174.600 120.200 ;
        RECT 175.800 117.900 176.200 120.200 ;
        RECT 179.800 117.900 180.200 120.200 ;
        RECT 181.400 117.900 181.800 120.200 ;
        RECT 183.000 117.900 183.400 120.200 ;
        RECT 184.600 117.900 185.000 120.200 ;
        RECT 169.400 115.900 169.800 116.200 ;
        RECT 171.000 115.900 171.500 116.000 ;
        RECT 186.200 115.900 186.600 120.200 ;
        RECT 189.000 117.900 189.400 120.200 ;
        RECT 190.600 117.900 191.000 120.200 ;
        RECT 193.400 116.000 193.800 120.200 ;
        RECT 195.800 116.000 196.200 120.200 ;
        RECT 198.600 117.900 199.000 120.200 ;
        RECT 200.200 117.900 200.600 120.200 ;
        RECT 203.000 115.900 203.400 120.200 ;
        RECT 135.500 115.600 149.000 115.900 ;
        RECT 169.400 115.600 182.900 115.900 ;
        RECT 135.500 115.500 135.900 115.600 ;
        RECT 182.500 115.500 182.900 115.600 ;
        RECT 1.400 100.800 1.800 105.100 ;
        RECT 4.200 100.800 4.600 103.100 ;
        RECT 5.800 100.800 6.200 103.100 ;
        RECT 8.600 100.800 9.000 105.000 ;
        RECT 10.200 100.800 10.600 103.100 ;
        RECT 11.800 100.800 12.200 105.100 ;
        RECT 13.900 100.800 14.300 103.100 ;
        RECT 15.000 100.800 15.400 103.100 ;
        RECT 16.600 100.800 17.000 103.100 ;
        RECT 18.000 100.800 18.400 105.100 ;
        RECT 20.600 100.800 21.000 104.900 ;
        RECT 22.200 100.800 22.600 103.100 ;
        RECT 23.800 100.800 24.200 105.100 ;
        RECT 25.900 100.800 26.300 103.100 ;
        RECT 27.000 100.800 27.400 103.100 ;
        RECT 29.400 100.800 29.800 104.500 ;
        RECT 32.100 100.800 32.500 103.100 ;
        RECT 34.200 100.800 34.600 105.100 ;
        RECT 35.000 100.800 35.400 103.100 ;
        RECT 36.600 100.800 37.000 105.100 ;
        RECT 38.700 100.800 39.100 103.100 ;
        RECT 41.400 100.800 41.800 104.500 ;
        RECT 43.800 100.800 44.200 104.500 ;
        RECT 46.200 100.800 46.600 105.100 ;
        RECT 47.800 100.800 48.200 104.500 ;
        RECT 51.800 100.800 52.200 104.500 ;
        RECT 53.400 100.800 53.800 105.100 ;
        RECT 54.200 100.800 54.600 105.100 ;
        RECT 55.800 100.800 56.200 104.500 ;
        RECT 57.400 100.800 57.800 105.100 ;
        RECT 60.600 100.800 61.000 105.100 ;
        RECT 61.400 100.800 61.800 105.100 ;
        RECT 63.000 100.800 63.400 104.500 ;
        RECT 64.600 100.800 65.000 103.100 ;
        RECT 67.800 100.800 68.200 104.500 ;
        RECT 69.400 100.800 69.800 105.100 ;
        RECT 72.600 100.800 73.000 105.100 ;
        RECT 73.400 100.800 73.800 105.100 ;
        RECT 76.600 100.800 77.000 105.000 ;
        RECT 79.400 100.800 79.800 103.100 ;
        RECT 81.000 100.800 81.400 103.100 ;
        RECT 83.800 100.800 84.200 105.100 ;
        RECT 85.400 100.800 85.800 103.100 ;
        RECT 87.000 100.800 87.400 103.100 ;
        RECT 89.400 100.800 89.800 105.100 ;
        RECT 90.500 100.800 90.900 103.100 ;
        RECT 92.600 100.800 93.000 105.100 ;
        RECT 93.400 100.800 93.800 105.100 ;
        RECT 95.000 100.800 95.400 104.500 ;
        RECT 97.400 100.800 97.800 103.100 ;
        RECT 98.200 100.800 98.600 103.100 ;
        RECT 99.800 100.800 100.200 103.100 ;
        RECT 102.500 100.800 102.900 103.100 ;
        RECT 104.600 100.800 105.000 105.100 ;
        RECT 106.200 100.800 106.600 105.100 ;
        RECT 109.000 100.800 109.400 103.100 ;
        RECT 110.600 100.800 111.000 103.100 ;
        RECT 113.400 100.800 113.800 105.000 ;
        RECT 115.800 100.800 116.200 104.500 ;
        RECT 117.400 100.800 117.800 105.100 ;
        RECT 119.000 100.800 119.400 105.000 ;
        RECT 121.800 100.800 122.200 103.100 ;
        RECT 123.400 100.800 123.800 103.100 ;
        RECT 126.200 100.800 126.600 105.100 ;
        RECT 127.800 100.800 128.200 105.100 ;
        RECT 131.800 100.800 132.200 104.500 ;
        RECT 134.200 100.800 134.600 104.900 ;
        RECT 136.800 100.800 137.200 105.100 ;
        RECT 139.000 100.800 139.400 103.100 ;
        RECT 140.600 100.800 141.000 105.100 ;
        RECT 143.400 100.800 143.800 103.100 ;
        RECT 145.000 100.800 145.400 103.100 ;
        RECT 147.800 100.800 148.200 105.000 ;
        RECT 151.800 100.800 152.200 105.000 ;
        RECT 154.600 100.800 155.000 103.100 ;
        RECT 156.200 100.800 156.600 103.100 ;
        RECT 159.000 100.800 159.400 105.100 ;
        RECT 161.400 100.800 161.800 104.500 ;
        RECT 165.400 100.800 165.800 105.100 ;
        RECT 167.000 100.800 167.400 104.500 ;
        RECT 170.200 100.800 170.600 104.500 ;
        RECT 171.800 100.800 172.200 105.100 ;
        RECT 172.900 100.800 173.300 103.100 ;
        RECT 175.000 100.800 175.400 105.100 ;
        RECT 176.600 100.800 177.000 103.100 ;
        RECT 178.200 100.800 178.600 105.100 ;
        RECT 181.000 100.800 181.400 103.100 ;
        RECT 182.600 100.800 183.000 103.100 ;
        RECT 185.400 100.800 185.800 105.000 ;
        RECT 187.800 100.800 188.200 104.900 ;
        RECT 190.400 100.800 190.800 105.100 ;
        RECT 192.600 100.800 193.000 104.900 ;
        RECT 195.200 100.800 195.600 105.100 ;
        RECT 196.600 100.800 197.000 105.100 ;
        RECT 198.700 100.800 199.100 103.100 ;
        RECT 199.800 100.800 200.200 103.100 ;
        RECT 201.400 100.800 201.800 103.100 ;
        RECT 202.200 100.800 202.600 103.100 ;
        RECT 203.800 100.800 204.200 103.100 ;
        RECT 0.200 100.200 205.400 100.800 ;
        RECT 0.600 95.900 1.000 100.200 ;
        RECT 2.200 95.900 2.600 100.200 ;
        RECT 3.800 95.900 4.200 100.200 ;
        RECT 5.400 95.900 5.800 100.200 ;
        RECT 7.000 95.900 7.400 100.200 ;
        RECT 8.600 96.000 9.000 100.200 ;
        RECT 11.400 97.900 11.800 100.200 ;
        RECT 13.000 97.900 13.400 100.200 ;
        RECT 15.800 95.900 16.200 100.200 ;
        RECT 17.400 95.900 17.800 100.200 ;
        RECT 19.500 97.900 19.900 100.200 ;
        RECT 20.600 97.900 21.000 100.200 ;
        RECT 22.200 97.900 22.600 100.200 ;
        RECT 23.800 96.500 24.200 100.200 ;
        RECT 26.200 97.900 26.600 100.200 ;
        RECT 28.600 96.500 29.000 100.200 ;
        RECT 31.800 96.500 32.200 100.200 ;
        RECT 34.200 95.900 34.600 100.200 ;
        RECT 36.300 97.900 36.700 100.200 ;
        RECT 37.400 95.900 37.800 100.200 ;
        RECT 39.500 97.900 39.900 100.200 ;
        RECT 42.200 96.500 42.600 100.200 ;
        RECT 44.100 97.900 44.500 100.200 ;
        RECT 46.200 95.900 46.600 100.200 ;
        RECT 47.000 95.900 47.400 100.200 ;
        RECT 50.200 95.900 50.600 100.200 ;
        RECT 52.600 95.900 53.000 100.200 ;
        RECT 54.200 96.500 54.600 100.200 ;
        RECT 56.100 97.900 56.500 100.200 ;
        RECT 58.200 95.900 58.600 100.200 ;
        RECT 59.800 96.500 60.200 100.200 ;
        RECT 63.800 96.500 64.200 100.200 ;
        RECT 66.200 96.500 66.600 100.200 ;
        RECT 67.800 95.900 68.200 100.200 ;
        RECT 68.600 95.900 69.000 100.200 ;
        RECT 70.200 95.900 70.600 100.200 ;
        RECT 71.800 95.900 72.200 100.200 ;
        RECT 72.600 95.900 73.000 100.200 ;
        RECT 75.800 95.900 76.200 100.200 ;
        RECT 76.900 97.900 77.300 100.200 ;
        RECT 79.000 95.900 79.400 100.200 ;
        RECT 80.100 97.900 80.500 100.200 ;
        RECT 82.200 95.900 82.600 100.200 ;
        RECT 83.300 97.900 83.700 100.200 ;
        RECT 85.400 95.900 85.800 100.200 ;
        RECT 86.200 95.900 86.600 100.200 ;
        RECT 89.400 95.900 89.800 100.200 ;
        RECT 91.800 96.500 92.200 100.200 ;
        RECT 93.700 97.900 94.100 100.200 ;
        RECT 95.800 95.900 96.200 100.200 ;
        RECT 96.600 95.900 97.000 100.200 ;
        RECT 98.200 96.500 98.600 100.200 ;
        RECT 99.800 95.900 100.200 100.200 ;
        RECT 101.400 96.500 101.800 100.200 ;
        RECT 105.400 96.000 105.800 100.200 ;
        RECT 108.200 97.900 108.600 100.200 ;
        RECT 109.800 97.900 110.200 100.200 ;
        RECT 112.600 95.900 113.000 100.200 ;
        RECT 114.200 95.900 114.600 100.200 ;
        RECT 116.300 97.900 116.700 100.200 ;
        RECT 117.400 97.900 117.800 100.200 ;
        RECT 119.000 97.900 119.400 100.200 ;
        RECT 120.100 97.900 120.500 100.200 ;
        RECT 122.200 95.900 122.600 100.200 ;
        RECT 123.000 95.900 123.400 100.200 ;
        RECT 124.600 96.500 125.000 100.200 ;
        RECT 127.000 96.500 127.400 100.200 ;
        RECT 128.600 95.900 129.000 100.200 ;
        RECT 130.200 96.000 130.600 100.200 ;
        RECT 133.000 97.900 133.400 100.200 ;
        RECT 134.600 97.900 135.000 100.200 ;
        RECT 137.400 95.900 137.800 100.200 ;
        RECT 139.800 96.500 140.200 100.200 ;
        RECT 143.800 95.900 144.200 100.200 ;
        RECT 144.600 95.900 145.000 100.200 ;
        RECT 146.700 97.900 147.100 100.200 ;
        RECT 148.600 96.500 149.000 100.200 ;
        RECT 151.800 96.500 152.200 100.200 ;
        RECT 153.400 95.900 153.800 100.200 ;
        RECT 156.900 95.900 157.300 100.200 ;
        RECT 160.600 96.500 161.000 100.200 ;
        RECT 162.200 97.900 162.600 100.200 ;
        RECT 163.800 97.900 164.200 100.200 ;
        RECT 164.900 97.900 165.300 100.200 ;
        RECT 167.000 95.900 167.400 100.200 ;
        RECT 168.100 97.900 168.500 100.200 ;
        RECT 170.200 95.900 170.600 100.200 ;
        RECT 171.000 95.900 171.400 100.200 ;
        RECT 173.100 97.900 173.500 100.200 ;
        RECT 175.800 96.500 176.200 100.200 ;
        RECT 178.200 96.100 178.600 100.200 ;
        RECT 180.800 95.900 181.200 100.200 ;
        RECT 183.000 97.900 183.400 100.200 ;
        RECT 184.600 95.900 185.000 100.200 ;
        RECT 187.400 97.900 187.800 100.200 ;
        RECT 189.000 97.900 189.400 100.200 ;
        RECT 191.800 96.000 192.200 100.200 ;
        RECT 194.200 97.900 194.600 100.200 ;
        RECT 195.800 95.900 196.200 100.200 ;
        RECT 198.600 97.900 199.000 100.200 ;
        RECT 200.200 97.900 200.600 100.200 ;
        RECT 203.000 96.000 203.400 100.200 ;
        RECT 1.400 80.800 1.800 85.100 ;
        RECT 4.200 80.800 4.600 83.100 ;
        RECT 5.800 80.800 6.200 83.100 ;
        RECT 8.600 80.800 9.000 85.000 ;
        RECT 10.200 80.800 10.600 83.100 ;
        RECT 11.800 80.800 12.200 83.100 ;
        RECT 12.900 80.800 13.300 83.100 ;
        RECT 15.000 80.800 15.400 85.100 ;
        RECT 15.800 80.800 16.200 83.100 ;
        RECT 17.400 80.800 17.800 83.100 ;
        RECT 19.000 80.800 19.400 84.500 ;
        RECT 21.700 80.800 22.100 83.100 ;
        RECT 23.800 80.800 24.200 85.100 ;
        RECT 25.400 80.800 25.800 85.000 ;
        RECT 28.200 80.800 28.600 83.100 ;
        RECT 29.800 80.800 30.200 83.100 ;
        RECT 32.600 80.800 33.000 85.100 ;
        RECT 34.200 80.800 34.600 85.100 ;
        RECT 38.200 80.800 38.600 84.500 ;
        RECT 40.600 80.800 41.000 84.500 ;
        RECT 43.300 80.800 43.700 83.100 ;
        RECT 45.400 80.800 45.800 85.100 ;
        RECT 47.000 80.800 47.400 83.100 ;
        RECT 50.200 80.800 50.600 85.100 ;
        RECT 53.000 80.800 53.400 83.100 ;
        RECT 54.600 80.800 55.000 83.100 ;
        RECT 57.400 80.800 57.800 85.000 ;
        RECT 59.000 80.800 59.400 83.100 ;
        RECT 60.600 80.800 61.000 83.100 ;
        RECT 61.700 80.800 62.100 83.100 ;
        RECT 63.800 80.800 64.200 85.100 ;
        RECT 65.400 80.800 65.800 84.500 ;
        RECT 67.000 80.800 67.400 85.100 ;
        RECT 68.100 80.800 68.500 83.100 ;
        RECT 70.200 80.800 70.600 85.100 ;
        RECT 71.300 80.800 71.700 83.100 ;
        RECT 73.400 80.800 73.800 85.100 ;
        RECT 75.800 80.800 76.200 84.500 ;
        RECT 77.400 80.800 77.800 85.100 ;
        RECT 79.000 80.800 79.400 84.500 ;
        RECT 80.600 80.800 81.000 85.100 ;
        RECT 82.700 80.800 83.100 83.100 ;
        RECT 84.100 80.800 84.500 83.100 ;
        RECT 86.200 80.800 86.600 85.100 ;
        RECT 87.000 80.800 87.400 85.100 ;
        RECT 88.600 80.800 89.000 85.100 ;
        RECT 90.200 80.800 90.600 85.100 ;
        RECT 91.800 80.800 92.200 84.500 ;
        RECT 94.500 80.800 94.900 83.100 ;
        RECT 96.600 80.800 97.000 85.100 ;
        RECT 98.200 80.800 98.600 83.100 ;
        RECT 99.000 80.800 99.400 83.100 ;
        RECT 100.600 80.800 101.000 83.100 ;
        RECT 103.300 80.800 103.700 83.100 ;
        RECT 105.400 80.800 105.800 85.100 ;
        RECT 107.000 80.800 107.400 85.100 ;
        RECT 109.800 80.800 110.200 83.100 ;
        RECT 111.400 80.800 111.800 83.100 ;
        RECT 114.200 80.800 114.600 85.000 ;
        RECT 117.400 80.800 117.800 84.500 ;
        RECT 119.800 80.800 120.200 85.100 ;
        RECT 122.600 80.800 123.000 83.100 ;
        RECT 124.200 80.800 124.600 83.100 ;
        RECT 127.000 80.800 127.400 85.000 ;
        RECT 128.600 80.800 129.000 85.100 ;
        RECT 132.600 80.800 133.000 84.500 ;
        RECT 135.000 80.800 135.400 84.500 ;
        RECT 136.600 80.800 137.000 85.100 ;
        RECT 138.200 80.800 138.600 85.100 ;
        RECT 141.000 80.800 141.400 83.100 ;
        RECT 142.600 80.800 143.000 83.100 ;
        RECT 145.400 80.800 145.800 85.000 ;
        RECT 147.300 80.800 147.700 83.100 ;
        RECT 149.400 80.800 149.800 85.100 ;
        RECT 151.000 80.800 151.400 84.900 ;
        RECT 153.600 80.800 154.000 85.100 ;
        RECT 158.200 80.800 158.600 84.500 ;
        RECT 160.600 80.800 161.000 83.100 ;
        RECT 162.200 80.800 162.600 85.100 ;
        RECT 165.000 80.800 165.400 83.100 ;
        RECT 166.600 80.800 167.000 83.100 ;
        RECT 169.400 80.800 169.800 85.000 ;
        RECT 171.000 80.800 171.400 85.100 ;
        RECT 173.100 80.800 173.500 83.100 ;
        RECT 174.200 80.800 174.600 83.100 ;
        RECT 175.800 80.800 176.200 83.100 ;
        RECT 176.900 80.800 177.300 83.100 ;
        RECT 179.000 80.800 179.400 85.100 ;
        RECT 180.600 80.800 181.000 85.100 ;
        RECT 183.400 80.800 183.800 83.100 ;
        RECT 185.000 80.800 185.400 83.100 ;
        RECT 187.800 80.800 188.200 85.000 ;
        RECT 190.000 80.800 190.400 85.100 ;
        RECT 192.600 80.800 193.000 84.900 ;
        RECT 195.000 80.800 195.400 83.100 ;
        RECT 196.600 80.800 197.000 85.100 ;
        RECT 199.400 80.800 199.800 83.100 ;
        RECT 201.000 80.800 201.400 83.100 ;
        RECT 203.800 80.800 204.200 85.000 ;
        RECT 0.200 80.200 205.400 80.800 ;
        RECT 1.400 76.000 1.800 80.200 ;
        RECT 4.200 77.900 4.600 80.200 ;
        RECT 5.800 77.900 6.200 80.200 ;
        RECT 8.600 75.900 9.000 80.200 ;
        RECT 10.200 75.900 10.600 80.200 ;
        RECT 14.200 76.500 14.600 80.200 ;
        RECT 16.100 77.900 16.500 80.200 ;
        RECT 18.200 75.900 18.600 80.200 ;
        RECT 19.800 76.000 20.200 80.200 ;
        RECT 22.600 77.900 23.000 80.200 ;
        RECT 24.200 77.900 24.600 80.200 ;
        RECT 27.000 75.900 27.400 80.200 ;
        RECT 28.600 77.900 29.000 80.200 ;
        RECT 30.200 77.900 30.600 80.200 ;
        RECT 31.800 77.900 32.200 80.200 ;
        RECT 33.400 76.000 33.800 80.200 ;
        RECT 36.200 77.900 36.600 80.200 ;
        RECT 37.800 77.900 38.200 80.200 ;
        RECT 40.600 75.900 41.000 80.200 ;
        RECT 42.200 77.900 42.600 80.200 ;
        RECT 43.800 77.900 44.200 80.200 ;
        RECT 44.900 77.900 45.300 80.200 ;
        RECT 47.000 75.900 47.400 80.200 ;
        RECT 47.800 75.900 48.200 80.200 ;
        RECT 49.900 77.900 50.300 80.200 ;
        RECT 52.600 75.900 53.000 80.200 ;
        RECT 54.700 77.900 55.100 80.200 ;
        RECT 55.800 75.900 56.200 80.200 ;
        RECT 57.400 76.500 57.800 80.200 ;
        RECT 60.600 75.900 61.000 80.200 ;
        RECT 61.400 75.900 61.800 80.200 ;
        RECT 64.600 75.900 65.000 80.200 ;
        RECT 65.400 75.900 65.800 80.200 ;
        RECT 67.500 77.900 67.900 80.200 ;
        RECT 68.600 75.900 69.000 80.200 ;
        RECT 70.700 77.900 71.100 80.200 ;
        RECT 71.800 75.900 72.200 80.200 ;
        RECT 75.000 75.900 75.400 80.200 ;
        RECT 75.800 75.900 76.200 80.200 ;
        RECT 79.000 75.900 79.400 80.200 ;
        RECT 79.800 75.900 80.200 80.200 ;
        RECT 83.000 75.900 83.400 80.200 ;
        RECT 83.800 75.900 84.200 80.200 ;
        RECT 85.900 77.900 86.300 80.200 ;
        RECT 88.600 76.500 89.000 80.200 ;
        RECT 90.200 75.900 90.600 80.200 ;
        RECT 93.400 75.900 93.800 80.200 ;
        RECT 94.200 75.900 94.600 80.200 ;
        RECT 97.400 75.900 97.800 80.200 ;
        RECT 100.200 77.900 100.600 80.200 ;
        RECT 101.800 77.900 102.200 80.200 ;
        RECT 104.600 76.000 105.000 80.200 ;
        RECT 107.800 77.900 108.200 80.200 ;
        RECT 109.400 77.900 109.800 80.200 ;
        RECT 110.500 77.900 110.900 80.200 ;
        RECT 112.600 75.900 113.000 80.200 ;
        RECT 113.400 75.900 113.800 80.200 ;
        RECT 116.100 77.900 116.500 80.200 ;
        RECT 118.200 75.900 118.600 80.200 ;
        RECT 119.800 75.900 120.200 80.200 ;
        RECT 122.600 77.900 123.000 80.200 ;
        RECT 124.200 77.900 124.600 80.200 ;
        RECT 127.000 76.000 127.400 80.200 ;
        RECT 128.600 75.900 129.000 80.200 ;
        RECT 131.000 75.900 131.400 80.200 ;
        RECT 135.000 76.500 135.400 80.200 ;
        RECT 136.600 75.900 137.000 80.200 ;
        RECT 138.700 77.900 139.100 80.200 ;
        RECT 139.800 77.900 140.200 80.200 ;
        RECT 141.400 77.900 141.800 80.200 ;
        RECT 143.000 76.000 143.400 80.200 ;
        RECT 145.800 77.900 146.200 80.200 ;
        RECT 147.400 77.900 147.800 80.200 ;
        RECT 150.200 75.900 150.600 80.200 ;
        RECT 154.200 76.500 154.600 80.200 ;
        RECT 156.600 77.900 157.000 80.200 ;
        RECT 158.500 77.900 158.900 80.200 ;
        RECT 160.600 75.900 161.000 80.200 ;
        RECT 161.400 77.900 161.800 80.200 ;
        RECT 163.000 77.900 163.400 80.200 ;
        RECT 163.800 75.900 164.200 80.200 ;
        RECT 167.800 76.500 168.200 80.200 ;
        RECT 170.200 76.500 170.600 80.200 ;
        RECT 171.800 75.900 172.200 80.200 ;
        RECT 174.200 76.500 174.600 80.200 ;
        RECT 175.800 75.900 176.200 80.200 ;
        RECT 179.800 76.500 180.200 80.200 ;
        RECT 182.200 75.900 182.600 80.200 ;
        RECT 185.000 77.900 185.400 80.200 ;
        RECT 186.600 77.900 187.000 80.200 ;
        RECT 189.400 76.000 189.800 80.200 ;
        RECT 191.800 77.900 192.200 80.200 ;
        RECT 193.400 76.500 193.800 80.200 ;
        RECT 196.600 75.900 197.000 80.200 ;
        RECT 199.400 77.900 199.800 80.200 ;
        RECT 201.000 77.900 201.400 80.200 ;
        RECT 203.800 76.000 204.200 80.200 ;
        RECT 1.400 60.800 1.800 65.000 ;
        RECT 4.200 60.800 4.600 63.100 ;
        RECT 5.800 60.800 6.200 63.100 ;
        RECT 8.600 60.800 9.000 65.100 ;
        RECT 10.500 60.800 10.900 63.100 ;
        RECT 12.600 60.800 13.000 65.100 ;
        RECT 13.400 60.800 13.800 63.100 ;
        RECT 15.000 60.800 15.400 63.100 ;
        RECT 16.600 60.800 17.000 65.000 ;
        RECT 19.400 60.800 19.800 63.100 ;
        RECT 21.000 60.800 21.400 63.100 ;
        RECT 23.800 60.800 24.200 65.100 ;
        RECT 25.400 60.800 25.800 65.100 ;
        RECT 27.500 60.800 27.900 63.100 ;
        RECT 28.600 60.800 29.000 65.100 ;
        RECT 30.700 60.800 31.100 63.100 ;
        RECT 31.800 60.800 32.200 63.100 ;
        RECT 33.400 60.800 33.800 63.100 ;
        RECT 35.000 60.800 35.400 65.000 ;
        RECT 37.800 60.800 38.200 63.100 ;
        RECT 39.400 60.800 39.800 63.100 ;
        RECT 42.200 60.800 42.600 65.100 ;
        RECT 43.800 60.800 44.200 65.100 ;
        RECT 45.900 60.800 46.300 63.100 ;
        RECT 47.800 60.800 48.200 64.500 ;
        RECT 51.800 60.800 52.200 65.100 ;
        RECT 53.900 60.800 54.300 63.100 ;
        RECT 55.300 60.800 55.700 63.100 ;
        RECT 57.400 60.800 57.800 65.100 ;
        RECT 58.200 60.800 58.600 63.100 ;
        RECT 59.800 60.800 60.200 63.100 ;
        RECT 61.400 60.800 61.800 65.000 ;
        RECT 64.200 60.800 64.600 63.100 ;
        RECT 65.800 60.800 66.200 63.100 ;
        RECT 68.600 60.800 69.000 65.100 ;
        RECT 71.000 60.800 71.400 64.500 ;
        RECT 73.400 60.800 73.800 65.100 ;
        RECT 76.600 60.800 77.000 64.500 ;
        RECT 78.200 60.800 78.600 65.100 ;
        RECT 79.000 60.800 79.400 63.100 ;
        RECT 80.600 60.800 81.000 63.100 ;
        RECT 81.700 60.800 82.100 63.100 ;
        RECT 83.800 60.800 84.200 65.100 ;
        RECT 84.900 60.800 85.300 63.100 ;
        RECT 87.000 60.800 87.400 65.100 ;
        RECT 87.800 60.800 88.200 63.100 ;
        RECT 89.400 60.800 89.800 63.100 ;
        RECT 90.500 60.800 90.900 63.100 ;
        RECT 92.600 60.800 93.000 65.100 ;
        RECT 93.400 60.800 93.800 63.100 ;
        RECT 95.000 60.800 95.400 63.100 ;
        RECT 96.100 60.800 96.500 63.100 ;
        RECT 98.200 60.800 98.600 65.100 ;
        RECT 100.600 60.800 101.000 64.500 ;
        RECT 104.100 60.800 104.500 63.100 ;
        RECT 106.200 60.800 106.600 65.100 ;
        RECT 107.800 60.800 108.200 65.000 ;
        RECT 110.600 60.800 111.000 63.100 ;
        RECT 112.200 60.800 112.600 63.100 ;
        RECT 115.000 60.800 115.400 65.100 ;
        RECT 117.400 60.800 117.800 64.500 ;
        RECT 120.600 60.800 121.000 65.100 ;
        RECT 123.400 60.800 123.800 63.100 ;
        RECT 125.000 60.800 125.400 63.100 ;
        RECT 127.800 60.800 128.200 65.000 ;
        RECT 131.000 60.800 131.400 64.500 ;
        RECT 132.600 60.800 133.000 63.100 ;
        RECT 134.200 60.800 134.600 63.100 ;
        RECT 135.300 60.800 135.700 63.100 ;
        RECT 137.400 60.800 137.800 65.100 ;
        RECT 139.000 60.800 139.400 64.500 ;
        RECT 142.200 60.800 142.600 64.500 ;
        RECT 143.800 60.800 144.200 65.100 ;
        RECT 144.900 60.800 145.300 63.100 ;
        RECT 147.000 60.800 147.400 65.100 ;
        RECT 148.600 60.800 149.000 64.500 ;
        RECT 151.000 60.800 151.400 65.100 ;
        RECT 153.100 60.800 153.500 63.100 ;
        RECT 156.600 60.800 157.000 65.000 ;
        RECT 159.400 60.800 159.800 63.100 ;
        RECT 161.000 60.800 161.400 63.100 ;
        RECT 163.800 60.800 164.200 65.100 ;
        RECT 166.200 60.800 166.600 64.900 ;
        RECT 168.800 60.800 169.200 65.100 ;
        RECT 171.000 60.800 171.400 63.100 ;
        RECT 172.600 60.800 173.000 65.100 ;
        RECT 175.400 60.800 175.800 63.100 ;
        RECT 177.000 60.800 177.400 63.100 ;
        RECT 179.800 60.800 180.200 65.000 ;
        RECT 182.000 60.800 182.400 65.100 ;
        RECT 184.600 60.800 185.000 64.900 ;
        RECT 187.000 60.800 187.400 64.500 ;
        RECT 189.700 60.800 190.100 63.100 ;
        RECT 191.800 60.800 192.200 65.100 ;
        RECT 192.600 60.800 193.000 65.100 ;
        RECT 194.200 60.800 194.600 65.100 ;
        RECT 195.300 60.800 195.700 63.100 ;
        RECT 197.400 60.800 197.800 65.100 ;
        RECT 198.200 60.800 198.600 65.100 ;
        RECT 202.200 60.800 202.600 64.500 ;
        RECT 0.200 60.200 205.400 60.800 ;
        RECT 1.400 56.000 1.800 60.200 ;
        RECT 4.200 57.900 4.600 60.200 ;
        RECT 5.800 57.900 6.200 60.200 ;
        RECT 8.600 55.900 9.000 60.200 ;
        RECT 11.000 56.000 11.400 60.200 ;
        RECT 13.800 57.900 14.200 60.200 ;
        RECT 15.400 57.900 15.800 60.200 ;
        RECT 18.200 55.900 18.600 60.200 ;
        RECT 19.800 55.900 20.200 60.200 ;
        RECT 21.900 57.900 22.300 60.200 ;
        RECT 23.000 57.900 23.400 60.200 ;
        RECT 24.600 57.900 25.000 60.200 ;
        RECT 26.200 56.000 26.600 60.200 ;
        RECT 29.000 57.900 29.400 60.200 ;
        RECT 30.600 57.900 31.000 60.200 ;
        RECT 33.400 55.900 33.800 60.200 ;
        RECT 35.000 57.900 35.400 60.200 ;
        RECT 36.600 57.900 37.000 60.200 ;
        RECT 37.700 57.900 38.100 60.200 ;
        RECT 39.800 55.900 40.200 60.200 ;
        RECT 40.600 55.900 41.000 60.200 ;
        RECT 42.700 57.900 43.100 60.200 ;
        RECT 44.600 56.000 45.000 60.200 ;
        RECT 47.400 57.900 47.800 60.200 ;
        RECT 49.000 57.900 49.400 60.200 ;
        RECT 51.800 55.900 52.200 60.200 ;
        RECT 55.000 55.900 55.400 60.200 ;
        RECT 57.100 57.900 57.500 60.200 ;
        RECT 58.200 57.900 58.600 60.200 ;
        RECT 59.800 57.900 60.200 60.200 ;
        RECT 60.900 57.900 61.300 60.200 ;
        RECT 63.000 55.900 63.400 60.200 ;
        RECT 64.600 56.500 65.000 60.200 ;
        RECT 67.800 56.000 68.200 60.200 ;
        RECT 70.600 57.900 71.000 60.200 ;
        RECT 72.200 57.900 72.600 60.200 ;
        RECT 75.000 55.900 75.400 60.200 ;
        RECT 76.600 55.900 77.000 60.200 ;
        RECT 78.700 57.900 79.100 60.200 ;
        RECT 79.800 57.900 80.200 60.200 ;
        RECT 81.400 57.900 81.800 60.200 ;
        RECT 83.800 56.500 84.200 60.200 ;
        RECT 85.700 57.900 86.100 60.200 ;
        RECT 87.800 55.900 88.200 60.200 ;
        RECT 88.600 55.900 89.000 60.200 ;
        RECT 90.700 57.900 91.100 60.200 ;
        RECT 91.800 57.900 92.200 60.200 ;
        RECT 93.400 57.900 93.800 60.200 ;
        RECT 95.000 56.000 95.400 60.200 ;
        RECT 97.800 57.900 98.200 60.200 ;
        RECT 99.400 57.900 99.800 60.200 ;
        RECT 102.200 55.900 102.600 60.200 ;
        RECT 105.700 57.900 106.100 60.200 ;
        RECT 107.800 55.900 108.200 60.200 ;
        RECT 109.400 57.900 109.800 60.200 ;
        RECT 110.200 57.900 110.600 60.200 ;
        RECT 111.800 57.900 112.200 60.200 ;
        RECT 112.900 57.900 113.300 60.200 ;
        RECT 115.000 55.900 115.400 60.200 ;
        RECT 116.600 56.500 117.000 60.200 ;
        RECT 119.800 55.900 120.200 60.200 ;
        RECT 122.600 57.900 123.000 60.200 ;
        RECT 124.200 57.900 124.600 60.200 ;
        RECT 127.000 56.000 127.400 60.200 ;
        RECT 128.600 55.900 129.000 60.200 ;
        RECT 130.700 57.900 131.100 60.200 ;
        RECT 131.800 57.900 132.200 60.200 ;
        RECT 133.400 57.900 133.800 60.200 ;
        RECT 135.000 56.000 135.400 60.200 ;
        RECT 137.800 57.900 138.200 60.200 ;
        RECT 139.400 57.900 139.800 60.200 ;
        RECT 142.200 55.900 142.600 60.200 ;
        RECT 144.600 56.500 145.000 60.200 ;
        RECT 146.200 55.900 146.600 60.200 ;
        RECT 147.800 55.900 148.200 60.200 ;
        RECT 150.600 57.900 151.000 60.200 ;
        RECT 152.200 57.900 152.600 60.200 ;
        RECT 155.000 56.000 155.400 60.200 ;
        RECT 159.000 57.900 159.400 60.200 ;
        RECT 160.600 55.900 161.000 60.200 ;
        RECT 163.400 57.900 163.800 60.200 ;
        RECT 165.000 57.900 165.400 60.200 ;
        RECT 167.800 56.000 168.200 60.200 ;
        RECT 170.200 56.100 170.600 60.200 ;
        RECT 172.800 55.900 173.200 60.200 ;
        RECT 175.000 56.500 175.400 60.200 ;
        RECT 177.700 57.900 178.100 60.200 ;
        RECT 179.800 55.900 180.200 60.200 ;
        RECT 181.400 56.000 181.800 60.200 ;
        RECT 184.200 57.900 184.600 60.200 ;
        RECT 185.800 57.900 186.200 60.200 ;
        RECT 188.600 55.900 189.000 60.200 ;
        RECT 190.200 57.900 190.600 60.200 ;
        RECT 191.800 57.900 192.200 60.200 ;
        RECT 193.400 57.900 193.800 60.200 ;
        RECT 195.000 56.500 195.400 60.200 ;
        RECT 199.000 55.900 199.400 60.200 ;
        RECT 199.800 57.900 200.200 60.200 ;
        RECT 201.400 57.900 201.800 60.200 ;
        RECT 203.800 56.500 204.200 60.200 ;
        RECT 0.600 40.800 1.000 45.100 ;
        RECT 2.200 40.800 2.600 45.100 ;
        RECT 3.800 40.800 4.200 45.100 ;
        RECT 5.400 40.800 5.800 45.100 ;
        RECT 7.000 40.800 7.400 45.100 ;
        RECT 7.800 40.800 8.200 45.100 ;
        RECT 11.800 40.800 12.200 44.500 ;
        RECT 13.400 40.800 13.800 43.100 ;
        RECT 15.000 40.800 15.400 43.100 ;
        RECT 16.100 40.800 16.500 43.100 ;
        RECT 18.200 40.800 18.600 45.100 ;
        RECT 19.000 40.800 19.400 45.100 ;
        RECT 21.100 40.800 21.500 43.100 ;
        RECT 22.200 40.800 22.600 43.100 ;
        RECT 23.800 40.800 24.200 43.100 ;
        RECT 25.400 40.800 25.800 45.000 ;
        RECT 28.200 40.800 28.600 43.100 ;
        RECT 29.800 40.800 30.200 43.100 ;
        RECT 32.600 40.800 33.000 45.100 ;
        RECT 34.200 40.800 34.600 45.100 ;
        RECT 36.300 40.800 36.700 43.100 ;
        RECT 37.400 40.800 37.800 43.100 ;
        RECT 39.000 40.800 39.400 43.100 ;
        RECT 40.600 40.800 41.000 45.000 ;
        RECT 43.400 40.800 43.800 43.100 ;
        RECT 45.000 40.800 45.400 43.100 ;
        RECT 47.800 40.800 48.200 45.100 ;
        RECT 51.000 40.800 51.400 45.100 ;
        RECT 53.100 40.800 53.500 43.100 ;
        RECT 54.200 40.800 54.600 45.100 ;
        RECT 56.300 40.800 56.700 43.100 ;
        RECT 58.200 40.800 58.600 44.500 ;
        RECT 59.800 40.800 60.200 45.100 ;
        RECT 61.400 40.800 61.800 45.000 ;
        RECT 64.200 40.800 64.600 43.100 ;
        RECT 65.800 40.800 66.200 43.100 ;
        RECT 68.600 40.800 69.000 45.100 ;
        RECT 71.000 40.800 71.400 45.000 ;
        RECT 73.800 40.800 74.200 43.100 ;
        RECT 75.400 40.800 75.800 43.100 ;
        RECT 78.200 40.800 78.600 45.100 ;
        RECT 79.800 40.800 80.200 43.100 ;
        RECT 82.000 40.800 82.400 45.100 ;
        RECT 84.600 40.800 85.000 44.900 ;
        RECT 87.800 40.800 88.200 45.100 ;
        RECT 89.400 40.800 89.800 44.500 ;
        RECT 91.800 40.800 92.200 45.100 ;
        RECT 93.900 40.800 94.300 43.100 ;
        RECT 95.300 40.800 95.700 43.100 ;
        RECT 97.400 40.800 97.800 45.100 ;
        RECT 99.000 40.800 99.400 44.500 ;
        RECT 100.600 40.800 101.000 45.100 ;
        RECT 103.800 40.800 104.200 44.500 ;
        RECT 107.000 40.800 107.400 44.500 ;
        RECT 111.000 40.800 111.400 44.500 ;
        RECT 112.900 40.800 113.300 43.100 ;
        RECT 115.000 40.800 115.400 45.100 ;
        RECT 117.400 40.800 117.800 45.100 ;
        RECT 119.000 40.800 119.400 45.100 ;
        RECT 121.800 40.800 122.200 43.100 ;
        RECT 123.400 40.800 123.800 43.100 ;
        RECT 126.200 40.800 126.600 45.000 ;
        RECT 128.100 40.800 128.500 43.100 ;
        RECT 130.200 40.800 130.600 45.100 ;
        RECT 131.000 40.800 131.400 45.100 ;
        RECT 132.600 40.800 133.000 44.500 ;
        RECT 135.000 40.800 135.400 45.100 ;
        RECT 137.800 40.800 138.200 43.100 ;
        RECT 139.400 40.800 139.800 43.100 ;
        RECT 142.200 40.800 142.600 45.000 ;
        RECT 143.800 40.800 144.200 45.100 ;
        RECT 147.800 40.800 148.200 44.500 ;
        RECT 149.700 40.800 150.100 43.100 ;
        RECT 151.800 40.800 152.200 45.100 ;
        RECT 154.200 40.800 154.600 45.100 ;
        RECT 155.800 40.800 156.200 45.100 ;
        RECT 157.400 40.800 157.800 44.900 ;
        RECT 160.000 40.800 160.400 45.100 ;
        RECT 162.200 40.800 162.600 44.500 ;
        RECT 164.900 40.800 165.300 43.100 ;
        RECT 167.000 40.800 167.400 45.100 ;
        RECT 167.800 40.800 168.200 43.100 ;
        RECT 169.400 40.800 169.800 43.100 ;
        RECT 170.200 40.800 170.600 43.100 ;
        RECT 171.800 40.800 172.200 43.100 ;
        RECT 172.600 40.800 173.000 45.100 ;
        RECT 174.200 40.800 174.600 45.100 ;
        RECT 175.800 40.800 176.200 45.000 ;
        RECT 178.600 40.800 179.000 43.100 ;
        RECT 180.200 40.800 180.600 43.100 ;
        RECT 183.000 40.800 183.400 45.100 ;
        RECT 184.600 40.800 185.000 43.100 ;
        RECT 187.000 40.800 187.400 44.900 ;
        RECT 189.600 40.800 190.000 45.100 ;
        RECT 191.800 40.800 192.200 45.000 ;
        RECT 194.600 40.800 195.000 43.100 ;
        RECT 196.200 40.800 196.600 43.100 ;
        RECT 199.000 40.800 199.400 45.100 ;
        RECT 200.600 40.800 201.000 45.100 ;
        RECT 202.200 40.800 202.600 45.100 ;
        RECT 203.000 40.800 203.400 45.100 ;
        RECT 0.200 40.200 205.400 40.800 ;
        RECT 0.600 37.900 1.000 40.200 ;
        RECT 3.000 36.000 3.400 40.200 ;
        RECT 5.800 37.900 6.200 40.200 ;
        RECT 7.400 37.900 7.800 40.200 ;
        RECT 10.200 35.900 10.600 40.200 ;
        RECT 12.400 35.900 12.800 40.200 ;
        RECT 15.000 36.100 15.400 40.200 ;
        RECT 16.600 37.900 17.000 40.200 ;
        RECT 19.000 36.100 19.400 40.200 ;
        RECT 21.600 35.900 22.000 40.200 ;
        RECT 23.800 36.000 24.200 40.200 ;
        RECT 26.600 37.900 27.000 40.200 ;
        RECT 28.200 37.900 28.600 40.200 ;
        RECT 31.000 35.900 31.400 40.200 ;
        RECT 32.600 35.900 33.000 40.200 ;
        RECT 34.700 37.900 35.100 40.200 ;
        RECT 35.800 37.900 36.200 40.200 ;
        RECT 37.400 37.900 37.800 40.200 ;
        RECT 38.200 37.900 38.600 40.200 ;
        RECT 40.600 36.500 41.000 40.200 ;
        RECT 43.000 35.900 43.400 40.200 ;
        RECT 45.100 37.900 45.500 40.200 ;
        RECT 47.000 36.500 47.400 40.200 ;
        RECT 51.800 36.500 52.200 40.200 ;
        RECT 54.200 35.900 54.600 40.200 ;
        RECT 56.600 35.900 57.000 40.200 ;
        RECT 59.300 37.900 59.700 40.200 ;
        RECT 61.400 35.900 61.800 40.200 ;
        RECT 62.200 35.900 62.600 40.200 ;
        RECT 63.800 36.500 64.200 40.200 ;
        RECT 65.400 35.900 65.800 40.200 ;
        RECT 67.500 37.900 67.900 40.200 ;
        RECT 68.600 37.900 69.000 40.200 ;
        RECT 70.200 37.900 70.600 40.200 ;
        RECT 71.000 35.900 71.400 40.200 ;
        RECT 72.600 36.500 73.000 40.200 ;
        RECT 74.200 35.900 74.600 40.200 ;
        RECT 75.800 35.900 76.200 40.200 ;
        RECT 77.400 35.900 77.800 40.200 ;
        RECT 78.200 35.900 78.600 40.200 ;
        RECT 80.900 37.900 81.300 40.200 ;
        RECT 83.000 35.900 83.400 40.200 ;
        RECT 83.800 35.900 84.200 40.200 ;
        RECT 85.900 37.900 86.300 40.200 ;
        RECT 87.000 37.900 87.400 40.200 ;
        RECT 88.600 37.900 89.000 40.200 ;
        RECT 90.200 35.900 90.600 40.200 ;
        RECT 93.000 37.900 93.400 40.200 ;
        RECT 94.600 37.900 95.000 40.200 ;
        RECT 97.400 36.000 97.800 40.200 ;
        RECT 100.600 35.900 101.000 40.200 ;
        RECT 103.000 35.900 103.400 40.200 ;
        RECT 106.200 35.900 106.600 40.200 ;
        RECT 107.600 35.900 108.000 40.200 ;
        RECT 110.200 36.100 110.600 40.200 ;
        RECT 112.600 36.500 113.000 40.200 ;
        RECT 115.800 37.900 116.200 40.200 ;
        RECT 117.400 35.900 117.800 40.200 ;
        RECT 120.200 37.900 120.600 40.200 ;
        RECT 121.800 37.900 122.200 40.200 ;
        RECT 124.600 36.000 125.000 40.200 ;
        RECT 126.200 35.900 126.600 40.200 ;
        RECT 130.200 36.500 130.600 40.200 ;
        RECT 132.400 35.900 132.800 40.200 ;
        RECT 135.000 36.100 135.400 40.200 ;
        RECT 137.400 37.900 137.800 40.200 ;
        RECT 139.000 35.900 139.400 40.200 ;
        RECT 141.800 37.900 142.200 40.200 ;
        RECT 143.400 37.900 143.800 40.200 ;
        RECT 146.200 36.000 146.600 40.200 ;
        RECT 147.800 35.900 148.200 40.200 ;
        RECT 149.400 35.900 149.800 40.200 ;
        RECT 151.000 35.900 151.400 40.200 ;
        RECT 152.600 35.900 153.000 40.200 ;
        RECT 154.200 35.900 154.600 40.200 ;
        RECT 157.400 37.900 157.800 40.200 ;
        RECT 159.000 35.900 159.400 40.200 ;
        RECT 161.800 37.900 162.200 40.200 ;
        RECT 163.400 37.900 163.800 40.200 ;
        RECT 166.200 36.000 166.600 40.200 ;
        RECT 167.800 35.900 168.200 40.200 ;
        RECT 171.800 36.500 172.200 40.200 ;
        RECT 174.200 36.100 174.600 40.200 ;
        RECT 176.800 35.900 177.200 40.200 ;
        RECT 179.000 37.900 179.400 40.200 ;
        RECT 179.800 35.900 180.200 40.200 ;
        RECT 183.800 36.500 184.200 40.200 ;
        RECT 186.200 35.900 186.600 40.200 ;
        RECT 189.000 37.900 189.400 40.200 ;
        RECT 190.600 37.900 191.000 40.200 ;
        RECT 193.400 36.000 193.800 40.200 ;
        RECT 195.800 35.900 196.200 40.200 ;
        RECT 198.600 37.900 199.000 40.200 ;
        RECT 200.200 37.900 200.600 40.200 ;
        RECT 203.000 36.000 203.400 40.200 ;
        RECT 1.400 20.800 1.800 25.100 ;
        RECT 4.200 20.800 4.600 23.100 ;
        RECT 5.800 20.800 6.200 23.100 ;
        RECT 8.600 20.800 9.000 25.000 ;
        RECT 11.000 20.800 11.400 25.100 ;
        RECT 13.800 20.800 14.200 23.100 ;
        RECT 15.400 20.800 15.800 23.100 ;
        RECT 18.200 20.800 18.600 25.000 ;
        RECT 20.600 20.800 21.000 25.000 ;
        RECT 23.400 20.800 23.800 23.100 ;
        RECT 25.000 20.800 25.400 23.100 ;
        RECT 27.800 20.800 28.200 25.100 ;
        RECT 29.400 20.800 29.800 23.100 ;
        RECT 31.000 20.800 31.400 23.100 ;
        RECT 32.100 20.800 32.500 23.100 ;
        RECT 34.200 20.800 34.600 25.100 ;
        RECT 35.800 20.800 36.200 25.000 ;
        RECT 38.600 20.800 39.000 23.100 ;
        RECT 40.200 20.800 40.600 23.100 ;
        RECT 43.000 20.800 43.400 25.100 ;
        RECT 44.600 20.800 45.000 25.100 ;
        RECT 46.700 20.800 47.100 23.100 ;
        RECT 47.800 20.800 48.200 23.100 ;
        RECT 49.400 20.800 49.800 23.100 ;
        RECT 51.800 20.800 52.200 25.100 ;
        RECT 53.400 20.800 53.800 24.500 ;
        RECT 55.000 20.800 55.400 25.100 ;
        RECT 57.100 20.800 57.500 23.100 ;
        RECT 59.800 20.800 60.200 24.500 ;
        RECT 61.400 20.800 61.800 25.100 ;
        RECT 64.100 20.800 64.500 23.100 ;
        RECT 66.200 20.800 66.600 25.100 ;
        RECT 67.000 20.800 67.400 25.100 ;
        RECT 69.100 20.800 69.500 23.100 ;
        RECT 70.500 20.800 70.900 23.100 ;
        RECT 72.600 20.800 73.000 25.100 ;
        RECT 74.000 20.800 74.400 25.100 ;
        RECT 76.600 20.800 77.000 24.900 ;
        RECT 78.200 20.800 78.600 23.100 ;
        RECT 79.800 20.800 80.200 23.100 ;
        RECT 80.900 20.800 81.300 23.100 ;
        RECT 83.000 20.800 83.400 25.100 ;
        RECT 83.800 20.800 84.200 25.100 ;
        RECT 85.900 20.800 86.300 23.100 ;
        RECT 87.800 20.800 88.200 24.900 ;
        RECT 90.400 20.800 90.800 25.100 ;
        RECT 91.800 20.800 92.200 25.100 ;
        RECT 93.900 20.800 94.300 23.100 ;
        RECT 95.000 20.800 95.400 25.100 ;
        RECT 97.100 20.800 97.500 23.100 ;
        RECT 99.000 20.800 99.400 24.900 ;
        RECT 101.600 20.800 102.000 25.100 ;
        RECT 106.200 20.800 106.600 24.500 ;
        RECT 107.800 20.800 108.200 25.100 ;
        RECT 111.800 20.800 112.200 24.500 ;
        RECT 113.700 20.800 114.100 23.100 ;
        RECT 115.800 20.800 116.200 25.100 ;
        RECT 116.900 20.800 117.300 23.100 ;
        RECT 119.000 20.800 119.400 25.100 ;
        RECT 120.100 20.800 120.500 23.100 ;
        RECT 122.200 20.800 122.600 25.100 ;
        RECT 123.000 20.800 123.400 25.100 ;
        RECT 125.100 20.800 125.500 23.100 ;
        RECT 127.000 20.800 127.400 24.500 ;
        RECT 129.700 20.800 130.100 23.100 ;
        RECT 131.800 20.800 132.200 25.100 ;
        RECT 133.400 20.800 133.800 25.100 ;
        RECT 136.200 20.800 136.600 23.100 ;
        RECT 137.800 20.800 138.200 23.100 ;
        RECT 140.600 20.800 141.000 25.000 ;
        RECT 142.200 20.800 142.600 25.100 ;
        RECT 145.400 20.800 145.800 25.100 ;
        RECT 148.200 20.800 148.600 23.100 ;
        RECT 149.800 20.800 150.200 23.100 ;
        RECT 152.600 20.800 153.000 25.000 ;
        RECT 156.600 20.800 157.000 24.500 ;
        RECT 159.000 20.800 159.400 25.100 ;
        RECT 163.000 20.800 163.400 24.500 ;
        RECT 164.900 20.800 165.300 23.100 ;
        RECT 167.000 20.800 167.400 25.100 ;
        RECT 168.600 20.800 169.000 25.100 ;
        RECT 171.400 20.800 171.800 23.100 ;
        RECT 173.000 20.800 173.400 23.100 ;
        RECT 175.800 20.800 176.200 25.000 ;
        RECT 178.200 20.800 178.600 25.100 ;
        RECT 181.000 20.800 181.400 23.100 ;
        RECT 182.600 20.800 183.000 23.100 ;
        RECT 185.400 20.800 185.800 25.000 ;
        RECT 187.800 20.800 188.200 24.900 ;
        RECT 190.400 20.800 190.800 25.100 ;
        RECT 192.600 20.800 193.000 25.100 ;
        RECT 194.200 20.800 194.600 23.100 ;
        RECT 195.800 20.800 196.200 24.900 ;
        RECT 198.400 20.800 198.800 25.100 ;
        RECT 200.600 20.800 201.000 24.500 ;
        RECT 203.000 20.800 203.400 24.500 ;
        RECT 0.200 20.200 205.400 20.800 ;
        RECT 1.400 16.000 1.800 20.200 ;
        RECT 4.200 17.900 4.600 20.200 ;
        RECT 5.800 17.900 6.200 20.200 ;
        RECT 8.600 15.900 9.000 20.200 ;
        RECT 11.000 16.500 11.400 20.200 ;
        RECT 15.000 15.900 15.400 20.200 ;
        RECT 16.600 16.000 17.000 20.200 ;
        RECT 19.400 17.900 19.800 20.200 ;
        RECT 21.000 17.900 21.400 20.200 ;
        RECT 23.800 15.900 24.200 20.200 ;
        RECT 25.400 15.900 25.800 20.200 ;
        RECT 27.500 17.900 27.900 20.200 ;
        RECT 28.600 17.900 29.000 20.200 ;
        RECT 30.200 17.900 30.600 20.200 ;
        RECT 31.000 15.900 31.400 20.200 ;
        RECT 33.100 17.900 33.500 20.200 ;
        RECT 34.200 17.900 34.600 20.200 ;
        RECT 35.800 17.900 36.200 20.200 ;
        RECT 36.600 17.900 37.000 20.200 ;
        RECT 38.200 17.900 38.600 20.200 ;
        RECT 39.800 17.900 40.200 20.200 ;
        RECT 41.400 16.000 41.800 20.200 ;
        RECT 44.200 17.900 44.600 20.200 ;
        RECT 45.800 17.900 46.200 20.200 ;
        RECT 48.600 15.900 49.000 20.200 ;
        RECT 51.800 15.900 52.200 20.200 ;
        RECT 53.900 17.900 54.300 20.200 ;
        RECT 55.000 17.900 55.400 20.200 ;
        RECT 56.600 17.900 57.000 20.200 ;
        RECT 57.400 15.900 57.800 20.200 ;
        RECT 61.400 15.900 61.800 20.200 ;
        RECT 63.000 15.900 63.400 20.200 ;
        RECT 65.800 17.900 66.200 20.200 ;
        RECT 67.400 17.900 67.800 20.200 ;
        RECT 70.200 16.000 70.600 20.200 ;
        RECT 71.800 15.900 72.200 20.200 ;
        RECT 73.900 17.900 74.300 20.200 ;
        RECT 75.000 15.900 75.400 20.200 ;
        RECT 77.100 17.900 77.500 20.200 ;
        RECT 78.200 15.900 78.600 20.200 ;
        RECT 81.400 15.900 81.800 20.200 ;
        RECT 82.200 17.900 82.600 20.200 ;
        RECT 83.800 17.900 84.200 20.200 ;
        RECT 85.400 17.900 85.800 20.200 ;
        RECT 86.500 17.900 86.900 20.200 ;
        RECT 88.600 15.900 89.000 20.200 ;
        RECT 90.200 16.000 90.600 20.200 ;
        RECT 93.000 17.900 93.400 20.200 ;
        RECT 94.600 17.900 95.000 20.200 ;
        RECT 97.400 15.900 97.800 20.200 ;
        RECT 99.800 17.900 100.200 20.200 ;
        RECT 100.600 15.900 101.000 20.200 ;
        RECT 105.400 15.900 105.800 20.200 ;
        RECT 108.200 17.900 108.600 20.200 ;
        RECT 109.800 17.900 110.200 20.200 ;
        RECT 112.600 16.000 113.000 20.200 ;
        RECT 114.200 17.900 114.600 20.200 ;
        RECT 115.800 17.900 116.200 20.200 ;
        RECT 116.900 17.900 117.300 20.200 ;
        RECT 119.000 15.900 119.400 20.200 ;
        RECT 120.600 16.000 121.000 20.200 ;
        RECT 123.400 17.900 123.800 20.200 ;
        RECT 125.000 17.900 125.400 20.200 ;
        RECT 127.800 15.900 128.200 20.200 ;
        RECT 129.400 15.900 129.800 20.200 ;
        RECT 131.000 15.900 131.400 20.200 ;
        RECT 132.600 15.900 133.000 20.200 ;
        RECT 134.200 15.900 134.600 20.200 ;
        RECT 135.800 15.900 136.200 20.200 ;
        RECT 137.400 16.100 137.800 20.200 ;
        RECT 140.000 15.900 140.400 20.200 ;
        RECT 141.400 15.900 141.800 20.200 ;
        RECT 145.400 16.500 145.800 20.200 ;
        RECT 147.800 15.900 148.200 20.200 ;
        RECT 150.600 17.900 151.000 20.200 ;
        RECT 152.200 17.900 152.600 20.200 ;
        RECT 155.000 16.000 155.400 20.200 ;
        RECT 158.200 15.900 158.600 20.200 ;
        RECT 162.200 16.500 162.600 20.200 ;
        RECT 163.800 15.900 164.200 20.200 ;
        RECT 167.800 16.500 168.200 20.200 ;
        RECT 169.400 15.900 169.800 20.200 ;
        RECT 171.000 15.900 171.400 20.200 ;
        RECT 172.600 15.900 173.000 20.200 ;
        RECT 174.200 15.900 174.600 20.200 ;
        RECT 175.800 15.900 176.200 20.200 ;
        RECT 176.600 15.900 177.000 20.200 ;
        RECT 180.600 16.500 181.000 20.200 ;
        RECT 182.200 15.900 182.600 20.200 ;
        RECT 186.200 16.500 186.600 20.200 ;
        RECT 188.600 16.000 189.000 20.200 ;
        RECT 191.400 17.900 191.800 20.200 ;
        RECT 193.000 17.900 193.400 20.200 ;
        RECT 195.800 15.900 196.200 20.200 ;
        RECT 198.200 16.500 198.600 20.200 ;
        RECT 200.600 17.900 201.000 20.200 ;
        RECT 202.200 16.500 202.600 20.200 ;
        RECT 0.600 0.800 1.000 5.100 ;
        RECT 2.200 0.800 2.600 5.100 ;
        RECT 3.800 0.800 4.200 5.100 ;
        RECT 5.400 0.800 5.800 5.100 ;
        RECT 7.000 0.800 7.400 5.100 ;
        RECT 7.800 0.800 8.200 5.100 ;
        RECT 9.400 0.800 9.800 5.100 ;
        RECT 11.000 0.800 11.400 5.100 ;
        RECT 12.600 0.800 13.000 5.100 ;
        RECT 14.200 0.800 14.600 5.100 ;
        RECT 15.800 0.800 16.200 5.000 ;
        RECT 18.600 0.800 19.000 3.100 ;
        RECT 20.200 0.800 20.600 3.100 ;
        RECT 23.000 0.800 23.400 5.100 ;
        RECT 24.600 0.800 25.000 5.100 ;
        RECT 28.600 0.800 29.000 4.500 ;
        RECT 31.000 0.800 31.400 5.000 ;
        RECT 33.800 0.800 34.200 3.100 ;
        RECT 35.400 0.800 35.800 3.100 ;
        RECT 38.200 0.800 38.600 5.100 ;
        RECT 40.100 0.800 40.500 3.100 ;
        RECT 42.200 0.800 42.600 5.100 ;
        RECT 43.800 0.800 44.200 5.100 ;
        RECT 46.600 0.800 47.000 3.100 ;
        RECT 48.200 0.800 48.600 3.100 ;
        RECT 51.000 0.800 51.400 5.000 ;
        RECT 55.000 0.800 55.400 5.000 ;
        RECT 57.800 0.800 58.200 3.100 ;
        RECT 59.400 0.800 59.800 3.100 ;
        RECT 62.200 0.800 62.600 5.100 ;
        RECT 63.800 0.800 64.200 3.100 ;
        RECT 65.400 0.800 65.800 3.100 ;
        RECT 66.500 0.800 66.900 3.100 ;
        RECT 68.600 0.800 69.000 5.100 ;
        RECT 70.200 0.800 70.600 5.000 ;
        RECT 73.000 0.800 73.400 3.100 ;
        RECT 74.600 0.800 75.000 3.100 ;
        RECT 77.400 0.800 77.800 5.100 ;
        RECT 79.000 0.800 79.400 3.100 ;
        RECT 80.600 0.800 81.000 3.100 ;
        RECT 82.200 0.800 82.600 5.100 ;
        RECT 85.000 0.800 85.400 3.100 ;
        RECT 86.600 0.800 87.000 3.100 ;
        RECT 89.400 0.800 89.800 5.000 ;
        RECT 91.800 0.800 92.200 5.100 ;
        RECT 94.600 0.800 95.000 3.100 ;
        RECT 96.200 0.800 96.600 3.100 ;
        RECT 99.000 0.800 99.400 5.000 ;
        RECT 103.000 0.800 103.400 5.100 ;
        RECT 105.800 0.800 106.200 3.100 ;
        RECT 107.400 0.800 107.800 3.100 ;
        RECT 110.200 0.800 110.600 5.000 ;
        RECT 111.800 0.800 112.200 3.100 ;
        RECT 113.400 0.800 113.800 3.100 ;
        RECT 114.500 0.800 114.900 3.100 ;
        RECT 116.600 0.800 117.000 5.100 ;
        RECT 119.000 0.800 119.400 5.100 ;
        RECT 121.400 0.800 121.800 4.500 ;
        RECT 123.800 0.800 124.200 5.100 ;
        RECT 126.600 0.800 127.000 3.100 ;
        RECT 128.200 0.800 128.600 3.100 ;
        RECT 131.000 0.800 131.400 5.000 ;
        RECT 133.400 0.800 133.800 3.100 ;
        RECT 135.000 0.800 135.400 5.100 ;
        RECT 137.800 0.800 138.200 3.100 ;
        RECT 139.400 0.800 139.800 3.100 ;
        RECT 142.200 0.800 142.600 5.000 ;
        RECT 143.800 0.800 144.200 5.100 ;
        RECT 145.400 0.800 145.800 5.100 ;
        RECT 147.000 0.800 147.400 5.100 ;
        RECT 148.600 0.800 149.000 5.100 ;
        RECT 150.200 0.800 150.600 5.100 ;
        RECT 153.400 0.800 153.800 5.100 ;
        RECT 156.200 0.800 156.600 3.100 ;
        RECT 157.800 0.800 158.200 3.100 ;
        RECT 160.600 0.800 161.000 5.000 ;
        RECT 162.200 0.800 162.600 3.100 ;
        RECT 164.600 0.800 165.000 5.100 ;
        RECT 167.400 0.800 167.800 3.100 ;
        RECT 169.000 0.800 169.400 3.100 ;
        RECT 171.800 0.800 172.200 5.000 ;
        RECT 174.200 0.800 174.600 5.100 ;
        RECT 177.000 0.800 177.400 3.100 ;
        RECT 178.600 0.800 179.000 3.100 ;
        RECT 181.400 0.800 181.800 5.000 ;
        RECT 183.800 0.800 184.200 5.100 ;
        RECT 186.600 0.800 187.000 3.100 ;
        RECT 188.200 0.800 188.600 3.100 ;
        RECT 191.000 0.800 191.400 5.000 ;
        RECT 193.400 0.800 193.800 5.000 ;
        RECT 196.200 0.800 196.600 3.100 ;
        RECT 197.800 0.800 198.200 3.100 ;
        RECT 200.600 0.800 201.000 5.100 ;
        RECT 202.200 0.800 202.600 5.100 ;
        RECT 203.800 0.800 204.200 5.100 ;
        RECT 0.200 0.200 205.400 0.800 ;
      LAYER via1 ;
        RECT 49.800 180.300 50.200 180.700 ;
        RECT 50.500 180.300 50.900 180.700 ;
        RECT 153.000 180.300 153.400 180.700 ;
        RECT 153.700 180.300 154.100 180.700 ;
        RECT 35.000 178.800 35.400 179.200 ;
        RECT 35.000 175.800 35.400 176.200 ;
        RECT 59.800 178.800 60.200 179.200 ;
        RECT 59.800 175.800 60.200 176.200 ;
        RECT 95.800 175.600 96.200 176.000 ;
        RECT 145.400 178.800 145.800 179.200 ;
        RECT 151.000 178.800 151.400 179.200 ;
        RECT 145.400 175.800 145.800 176.200 ;
        RECT 151.000 175.800 151.400 176.200 ;
        RECT 175.800 178.800 176.200 179.200 ;
        RECT 175.800 175.800 176.200 176.200 ;
        RECT 31.800 165.000 32.200 165.400 ;
        RECT 49.400 165.000 49.800 165.400 ;
        RECT 15.800 161.800 16.200 162.200 ;
        RECT 31.800 161.800 32.200 162.200 ;
        RECT 49.400 162.700 49.800 163.100 ;
        RECT 150.200 161.800 150.600 162.200 ;
        RECT 167.000 161.800 167.400 162.200 ;
        RECT 49.800 160.300 50.200 160.700 ;
        RECT 50.500 160.300 50.900 160.700 ;
        RECT 153.000 160.300 153.400 160.700 ;
        RECT 153.700 160.300 154.100 160.700 ;
        RECT 32.600 158.800 33.000 159.200 ;
        RECT 32.600 155.800 33.000 156.200 ;
        RECT 79.800 158.800 80.200 159.200 ;
        RECT 79.800 155.800 80.200 156.200 ;
        RECT 139.800 158.800 140.200 159.200 ;
        RECT 157.400 158.800 157.800 159.200 ;
        RECT 163.000 158.800 163.400 159.200 ;
        RECT 139.800 155.800 140.200 156.200 ;
        RECT 157.400 155.800 157.800 156.200 ;
        RECT 163.000 155.800 163.400 156.200 ;
        RECT 80.600 145.000 81.000 145.400 ;
        RECT 80.600 141.800 81.000 142.200 ;
        RECT 49.800 140.300 50.200 140.700 ;
        RECT 50.500 140.300 50.900 140.700 ;
        RECT 153.000 140.300 153.400 140.700 ;
        RECT 153.700 140.300 154.100 140.700 ;
        RECT 15.800 138.800 16.200 139.200 ;
        RECT 35.800 138.800 36.200 139.200 ;
        RECT 15.800 135.800 16.200 136.200 ;
        RECT 35.800 135.800 36.200 136.200 ;
        RECT 49.800 120.300 50.200 120.700 ;
        RECT 50.500 120.300 50.900 120.700 ;
        RECT 153.000 120.300 153.400 120.700 ;
        RECT 153.700 120.300 154.100 120.700 ;
        RECT 147.000 115.600 147.400 116.000 ;
        RECT 171.000 115.600 171.400 116.000 ;
        RECT 49.800 100.300 50.200 100.700 ;
        RECT 50.500 100.300 50.900 100.700 ;
        RECT 153.000 100.300 153.400 100.700 ;
        RECT 153.700 100.300 154.100 100.700 ;
        RECT 49.800 80.300 50.200 80.700 ;
        RECT 50.500 80.300 50.900 80.700 ;
        RECT 153.000 80.300 153.400 80.700 ;
        RECT 153.700 80.300 154.100 80.700 ;
        RECT 49.800 60.300 50.200 60.700 ;
        RECT 50.500 60.300 50.900 60.700 ;
        RECT 153.000 60.300 153.400 60.700 ;
        RECT 153.700 60.300 154.100 60.700 ;
        RECT 49.800 40.300 50.200 40.700 ;
        RECT 50.500 40.300 50.900 40.700 ;
        RECT 153.000 40.300 153.400 40.700 ;
        RECT 153.700 40.300 154.100 40.700 ;
        RECT 49.800 20.300 50.200 20.700 ;
        RECT 50.500 20.300 50.900 20.700 ;
        RECT 153.000 20.300 153.400 20.700 ;
        RECT 153.700 20.300 154.100 20.700 ;
        RECT 49.800 0.300 50.200 0.700 ;
        RECT 50.500 0.300 50.900 0.700 ;
        RECT 153.000 0.300 153.400 0.700 ;
        RECT 153.700 0.300 154.100 0.700 ;
      LAYER metal2 ;
        RECT 49.600 180.300 51.200 180.700 ;
        RECT 152.800 180.300 154.400 180.700 ;
        RECT 35.000 178.800 35.400 179.200 ;
        RECT 59.800 178.800 60.200 179.200 ;
        RECT 145.400 178.800 145.800 179.200 ;
        RECT 151.000 178.800 151.400 179.200 ;
        RECT 175.800 178.800 176.200 179.200 ;
        RECT 35.000 176.200 35.300 178.800 ;
        RECT 59.800 176.200 60.100 178.800 ;
        RECT 95.800 177.900 96.200 178.300 ;
        RECT 35.000 175.800 35.400 176.200 ;
        RECT 59.800 175.800 60.200 176.200 ;
        RECT 95.800 176.000 96.100 177.900 ;
        RECT 145.400 176.200 145.700 178.800 ;
        RECT 151.000 176.200 151.300 178.800 ;
        RECT 175.800 176.200 176.100 178.800 ;
        RECT 95.800 175.600 96.200 176.000 ;
        RECT 145.400 175.800 145.800 176.200 ;
        RECT 151.000 175.800 151.400 176.200 ;
        RECT 175.800 175.800 176.200 176.200 ;
        RECT 15.800 164.800 16.200 165.200 ;
        RECT 31.800 165.000 32.200 165.400 ;
        RECT 49.400 165.000 49.800 165.400 ;
        RECT 15.800 162.200 16.100 164.800 ;
        RECT 31.800 162.200 32.100 165.000 ;
        RECT 49.400 163.100 49.700 165.000 ;
        RECT 150.200 164.800 150.600 165.200 ;
        RECT 167.000 164.800 167.400 165.200 ;
        RECT 49.400 162.700 49.800 163.100 ;
        RECT 150.200 162.200 150.500 164.800 ;
        RECT 167.000 162.200 167.300 164.800 ;
        RECT 15.800 161.800 16.200 162.200 ;
        RECT 31.800 161.800 32.200 162.200 ;
        RECT 150.200 161.800 150.600 162.200 ;
        RECT 167.000 161.800 167.400 162.200 ;
        RECT 49.600 160.300 51.200 160.700 ;
        RECT 152.800 160.300 154.400 160.700 ;
        RECT 32.600 158.800 33.000 159.200 ;
        RECT 79.800 158.800 80.200 159.200 ;
        RECT 139.800 158.800 140.200 159.200 ;
        RECT 157.400 158.800 157.800 159.200 ;
        RECT 163.000 158.800 163.400 159.200 ;
        RECT 32.600 156.200 32.900 158.800 ;
        RECT 79.800 156.200 80.100 158.800 ;
        RECT 139.800 156.200 140.100 158.800 ;
        RECT 157.400 156.200 157.700 158.800 ;
        RECT 163.000 156.200 163.300 158.800 ;
        RECT 32.600 155.800 33.000 156.200 ;
        RECT 79.800 155.800 80.200 156.200 ;
        RECT 139.800 155.800 140.200 156.200 ;
        RECT 157.400 155.800 157.800 156.200 ;
        RECT 163.000 155.800 163.400 156.200 ;
        RECT 80.600 145.000 81.000 145.400 ;
        RECT 80.600 142.200 80.900 145.000 ;
        RECT 80.600 141.800 81.000 142.200 ;
        RECT 49.600 140.300 51.200 140.700 ;
        RECT 152.800 140.300 154.400 140.700 ;
        RECT 15.800 138.800 16.200 139.200 ;
        RECT 35.800 138.800 36.200 139.200 ;
        RECT 15.800 136.200 16.100 138.800 ;
        RECT 35.800 136.200 36.100 138.800 ;
        RECT 15.800 135.800 16.200 136.200 ;
        RECT 35.800 135.800 36.200 136.200 ;
        RECT 49.600 120.300 51.200 120.700 ;
        RECT 152.800 120.300 154.400 120.700 ;
        RECT 147.000 117.900 147.400 118.300 ;
        RECT 171.000 117.900 171.400 118.300 ;
        RECT 147.000 116.000 147.300 117.900 ;
        RECT 171.000 116.000 171.300 117.900 ;
        RECT 147.000 115.600 147.400 116.000 ;
        RECT 171.000 115.600 171.400 116.000 ;
        RECT 49.600 100.300 51.200 100.700 ;
        RECT 152.800 100.300 154.400 100.700 ;
        RECT 49.600 80.300 51.200 80.700 ;
        RECT 152.800 80.300 154.400 80.700 ;
        RECT 49.600 60.300 51.200 60.700 ;
        RECT 152.800 60.300 154.400 60.700 ;
        RECT 49.600 40.300 51.200 40.700 ;
        RECT 152.800 40.300 154.400 40.700 ;
        RECT 49.600 20.300 51.200 20.700 ;
        RECT 152.800 20.300 154.400 20.700 ;
        RECT 49.600 0.300 51.200 0.700 ;
        RECT 152.800 0.300 154.400 0.700 ;
      LAYER via2 ;
        RECT 49.800 180.300 50.200 180.700 ;
        RECT 50.500 180.300 50.900 180.700 ;
        RECT 153.000 180.300 153.400 180.700 ;
        RECT 153.700 180.300 154.100 180.700 ;
        RECT 49.800 160.300 50.200 160.700 ;
        RECT 50.500 160.300 50.900 160.700 ;
        RECT 153.000 160.300 153.400 160.700 ;
        RECT 153.700 160.300 154.100 160.700 ;
        RECT 49.800 140.300 50.200 140.700 ;
        RECT 50.500 140.300 50.900 140.700 ;
        RECT 153.000 140.300 153.400 140.700 ;
        RECT 153.700 140.300 154.100 140.700 ;
        RECT 49.800 120.300 50.200 120.700 ;
        RECT 50.500 120.300 50.900 120.700 ;
        RECT 153.000 120.300 153.400 120.700 ;
        RECT 153.700 120.300 154.100 120.700 ;
        RECT 49.800 100.300 50.200 100.700 ;
        RECT 50.500 100.300 50.900 100.700 ;
        RECT 153.000 100.300 153.400 100.700 ;
        RECT 153.700 100.300 154.100 100.700 ;
        RECT 49.800 80.300 50.200 80.700 ;
        RECT 50.500 80.300 50.900 80.700 ;
        RECT 153.000 80.300 153.400 80.700 ;
        RECT 153.700 80.300 154.100 80.700 ;
        RECT 49.800 60.300 50.200 60.700 ;
        RECT 50.500 60.300 50.900 60.700 ;
        RECT 153.000 60.300 153.400 60.700 ;
        RECT 153.700 60.300 154.100 60.700 ;
        RECT 49.800 40.300 50.200 40.700 ;
        RECT 50.500 40.300 50.900 40.700 ;
        RECT 153.000 40.300 153.400 40.700 ;
        RECT 153.700 40.300 154.100 40.700 ;
        RECT 49.800 20.300 50.200 20.700 ;
        RECT 50.500 20.300 50.900 20.700 ;
        RECT 153.000 20.300 153.400 20.700 ;
        RECT 153.700 20.300 154.100 20.700 ;
        RECT 49.800 0.300 50.200 0.700 ;
        RECT 50.500 0.300 50.900 0.700 ;
        RECT 153.000 0.300 153.400 0.700 ;
        RECT 153.700 0.300 154.100 0.700 ;
      LAYER metal3 ;
        RECT 49.600 180.300 51.200 180.700 ;
        RECT 152.800 180.300 154.400 180.700 ;
        RECT 49.600 160.300 51.200 160.700 ;
        RECT 152.800 160.300 154.400 160.700 ;
        RECT 49.600 140.300 51.200 140.700 ;
        RECT 152.800 140.300 154.400 140.700 ;
        RECT 49.600 120.300 51.200 120.700 ;
        RECT 152.800 120.300 154.400 120.700 ;
        RECT 49.600 100.300 51.200 100.700 ;
        RECT 152.800 100.300 154.400 100.700 ;
        RECT 49.600 80.300 51.200 80.700 ;
        RECT 152.800 80.300 154.400 80.700 ;
        RECT 49.600 60.300 51.200 60.700 ;
        RECT 152.800 60.300 154.400 60.700 ;
        RECT 49.600 40.300 51.200 40.700 ;
        RECT 152.800 40.300 154.400 40.700 ;
        RECT 49.600 20.300 51.200 20.700 ;
        RECT 152.800 20.300 154.400 20.700 ;
        RECT 49.600 0.300 51.200 0.700 ;
        RECT 152.800 0.300 154.400 0.700 ;
      LAYER via3 ;
        RECT 49.800 180.300 50.200 180.700 ;
        RECT 50.600 180.300 51.000 180.700 ;
        RECT 153.000 180.300 153.400 180.700 ;
        RECT 153.800 180.300 154.200 180.700 ;
        RECT 49.800 160.300 50.200 160.700 ;
        RECT 50.600 160.300 51.000 160.700 ;
        RECT 153.000 160.300 153.400 160.700 ;
        RECT 153.800 160.300 154.200 160.700 ;
        RECT 49.800 140.300 50.200 140.700 ;
        RECT 50.600 140.300 51.000 140.700 ;
        RECT 153.000 140.300 153.400 140.700 ;
        RECT 153.800 140.300 154.200 140.700 ;
        RECT 49.800 120.300 50.200 120.700 ;
        RECT 50.600 120.300 51.000 120.700 ;
        RECT 153.000 120.300 153.400 120.700 ;
        RECT 153.800 120.300 154.200 120.700 ;
        RECT 49.800 100.300 50.200 100.700 ;
        RECT 50.600 100.300 51.000 100.700 ;
        RECT 153.000 100.300 153.400 100.700 ;
        RECT 153.800 100.300 154.200 100.700 ;
        RECT 49.800 80.300 50.200 80.700 ;
        RECT 50.600 80.300 51.000 80.700 ;
        RECT 153.000 80.300 153.400 80.700 ;
        RECT 153.800 80.300 154.200 80.700 ;
        RECT 49.800 60.300 50.200 60.700 ;
        RECT 50.600 60.300 51.000 60.700 ;
        RECT 153.000 60.300 153.400 60.700 ;
        RECT 153.800 60.300 154.200 60.700 ;
        RECT 49.800 40.300 50.200 40.700 ;
        RECT 50.600 40.300 51.000 40.700 ;
        RECT 153.000 40.300 153.400 40.700 ;
        RECT 153.800 40.300 154.200 40.700 ;
        RECT 49.800 20.300 50.200 20.700 ;
        RECT 50.600 20.300 51.000 20.700 ;
        RECT 153.000 20.300 153.400 20.700 ;
        RECT 153.800 20.300 154.200 20.700 ;
        RECT 49.800 0.300 50.200 0.700 ;
        RECT 50.600 0.300 51.000 0.700 ;
        RECT 153.000 0.300 153.400 0.700 ;
        RECT 153.800 0.300 154.200 0.700 ;
      LAYER metal4 ;
        RECT 49.600 180.300 51.200 180.700 ;
        RECT 152.800 180.300 154.400 180.700 ;
        RECT 49.600 160.300 51.200 160.700 ;
        RECT 152.800 160.300 154.400 160.700 ;
        RECT 49.600 140.300 51.200 140.700 ;
        RECT 152.800 140.300 154.400 140.700 ;
        RECT 49.600 120.300 51.200 120.700 ;
        RECT 152.800 120.300 154.400 120.700 ;
        RECT 49.600 100.300 51.200 100.700 ;
        RECT 152.800 100.300 154.400 100.700 ;
        RECT 49.600 80.300 51.200 80.700 ;
        RECT 152.800 80.300 154.400 80.700 ;
        RECT 49.600 60.300 51.200 60.700 ;
        RECT 152.800 60.300 154.400 60.700 ;
        RECT 49.600 40.300 51.200 40.700 ;
        RECT 152.800 40.300 154.400 40.700 ;
        RECT 49.600 20.300 51.200 20.700 ;
        RECT 152.800 20.300 154.400 20.700 ;
        RECT 49.600 0.300 51.200 0.700 ;
        RECT 152.800 0.300 154.400 0.700 ;
      LAYER via4 ;
        RECT 49.800 180.300 50.200 180.700 ;
        RECT 50.500 180.300 50.900 180.700 ;
        RECT 153.000 180.300 153.400 180.700 ;
        RECT 153.700 180.300 154.100 180.700 ;
        RECT 49.800 160.300 50.200 160.700 ;
        RECT 50.500 160.300 50.900 160.700 ;
        RECT 153.000 160.300 153.400 160.700 ;
        RECT 153.700 160.300 154.100 160.700 ;
        RECT 49.800 140.300 50.200 140.700 ;
        RECT 50.500 140.300 50.900 140.700 ;
        RECT 153.000 140.300 153.400 140.700 ;
        RECT 153.700 140.300 154.100 140.700 ;
        RECT 49.800 120.300 50.200 120.700 ;
        RECT 50.500 120.300 50.900 120.700 ;
        RECT 153.000 120.300 153.400 120.700 ;
        RECT 153.700 120.300 154.100 120.700 ;
        RECT 49.800 100.300 50.200 100.700 ;
        RECT 50.500 100.300 50.900 100.700 ;
        RECT 153.000 100.300 153.400 100.700 ;
        RECT 153.700 100.300 154.100 100.700 ;
        RECT 49.800 80.300 50.200 80.700 ;
        RECT 50.500 80.300 50.900 80.700 ;
        RECT 153.000 80.300 153.400 80.700 ;
        RECT 153.700 80.300 154.100 80.700 ;
        RECT 49.800 60.300 50.200 60.700 ;
        RECT 50.500 60.300 50.900 60.700 ;
        RECT 153.000 60.300 153.400 60.700 ;
        RECT 153.700 60.300 154.100 60.700 ;
        RECT 49.800 40.300 50.200 40.700 ;
        RECT 50.500 40.300 50.900 40.700 ;
        RECT 153.000 40.300 153.400 40.700 ;
        RECT 153.700 40.300 154.100 40.700 ;
        RECT 49.800 20.300 50.200 20.700 ;
        RECT 50.500 20.300 50.900 20.700 ;
        RECT 153.000 20.300 153.400 20.700 ;
        RECT 153.700 20.300 154.100 20.700 ;
        RECT 49.800 0.300 50.200 0.700 ;
        RECT 50.500 0.300 50.900 0.700 ;
        RECT 153.000 0.300 153.400 0.700 ;
        RECT 153.700 0.300 154.100 0.700 ;
      LAYER metal5 ;
        RECT 49.600 180.200 51.200 180.700 ;
        RECT 152.800 180.200 154.400 180.700 ;
        RECT 49.600 160.200 51.200 160.700 ;
        RECT 152.800 160.200 154.400 160.700 ;
        RECT 49.600 140.200 51.200 140.700 ;
        RECT 152.800 140.200 154.400 140.700 ;
        RECT 49.600 120.200 51.200 120.700 ;
        RECT 152.800 120.200 154.400 120.700 ;
        RECT 49.600 100.200 51.200 100.700 ;
        RECT 152.800 100.200 154.400 100.700 ;
        RECT 49.600 80.200 51.200 80.700 ;
        RECT 152.800 80.200 154.400 80.700 ;
        RECT 49.600 60.200 51.200 60.700 ;
        RECT 152.800 60.200 154.400 60.700 ;
        RECT 49.600 40.200 51.200 40.700 ;
        RECT 152.800 40.200 154.400 40.700 ;
        RECT 49.600 20.200 51.200 20.700 ;
        RECT 152.800 20.200 154.400 20.700 ;
        RECT 49.600 0.200 51.200 0.700 ;
        RECT 152.800 0.200 154.400 0.700 ;
      LAYER via5 ;
        RECT 50.600 180.200 51.100 180.700 ;
        RECT 153.800 180.200 154.300 180.700 ;
        RECT 50.600 160.200 51.100 160.700 ;
        RECT 153.800 160.200 154.300 160.700 ;
        RECT 50.600 140.200 51.100 140.700 ;
        RECT 153.800 140.200 154.300 140.700 ;
        RECT 50.600 120.200 51.100 120.700 ;
        RECT 153.800 120.200 154.300 120.700 ;
        RECT 50.600 100.200 51.100 100.700 ;
        RECT 153.800 100.200 154.300 100.700 ;
        RECT 50.600 80.200 51.100 80.700 ;
        RECT 153.800 80.200 154.300 80.700 ;
        RECT 50.600 60.200 51.100 60.700 ;
        RECT 153.800 60.200 154.300 60.700 ;
        RECT 50.600 40.200 51.100 40.700 ;
        RECT 153.800 40.200 154.300 40.700 ;
        RECT 50.600 20.200 51.100 20.700 ;
        RECT 153.800 20.200 154.300 20.700 ;
        RECT 50.600 0.200 51.100 0.700 ;
        RECT 153.800 0.200 154.300 0.700 ;
      LAYER metal6 ;
        RECT 49.600 -3.000 51.200 183.000 ;
        RECT 152.800 -3.000 154.400 183.000 ;
    END
  END vdd
  PIN gnd
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 1.400 170.800 1.800 173.100 ;
        RECT 3.800 170.800 4.200 173.100 ;
        RECT 5.400 170.800 5.800 173.100 ;
        RECT 7.000 170.800 7.400 173.100 ;
        RECT 8.600 170.800 9.000 173.100 ;
        RECT 10.200 170.800 10.600 173.100 ;
        RECT 11.800 170.800 12.200 173.100 ;
        RECT 13.400 170.800 13.800 173.100 ;
        RECT 15.800 170.800 16.200 173.100 ;
        RECT 18.200 170.800 18.600 173.100 ;
        RECT 19.800 170.800 20.200 172.100 ;
        RECT 23.000 170.800 23.400 173.100 ;
        RECT 28.600 170.800 29.000 172.100 ;
        RECT 30.200 170.800 30.600 172.100 ;
        RECT 35.000 170.800 35.400 173.100 ;
        RECT 37.400 170.800 37.800 173.100 ;
        RECT 39.000 170.800 39.400 173.100 ;
        RECT 41.400 170.800 41.800 173.100 ;
        RECT 44.600 170.800 45.000 172.100 ;
        RECT 47.800 170.800 48.200 173.100 ;
        RECT 53.400 170.800 53.800 172.100 ;
        RECT 55.000 170.800 55.400 172.100 ;
        RECT 59.800 170.800 60.200 173.100 ;
        RECT 63.000 170.800 63.400 173.000 ;
        RECT 65.800 170.800 66.200 172.100 ;
        RECT 67.400 170.800 67.900 172.100 ;
        RECT 70.200 170.800 70.600 173.100 ;
        RECT 72.600 170.800 73.000 173.000 ;
        RECT 75.400 170.800 75.800 172.100 ;
        RECT 77.000 170.800 77.500 172.100 ;
        RECT 79.800 170.800 80.200 173.100 ;
        RECT 81.400 170.800 81.800 173.100 ;
        RECT 83.000 170.800 83.400 173.100 ;
        RECT 84.600 170.800 85.000 173.100 ;
        RECT 85.400 170.800 85.800 173.100 ;
        RECT 87.000 170.800 87.400 173.100 ;
        RECT 88.600 170.800 89.000 173.100 ;
        RECT 90.200 170.800 90.600 173.100 ;
        RECT 91.800 170.800 92.200 173.100 ;
        RECT 94.200 170.800 94.600 173.100 ;
        RECT 99.000 170.800 99.400 172.100 ;
        RECT 100.600 170.800 101.000 172.100 ;
        RECT 106.200 170.800 106.600 173.100 ;
        RECT 109.400 170.800 109.800 172.100 ;
        RECT 112.600 170.800 113.000 173.100 ;
        RECT 114.200 170.800 114.600 173.100 ;
        RECT 115.000 170.800 115.400 173.100 ;
        RECT 116.600 170.800 117.000 173.100 ;
        RECT 118.200 170.800 118.600 173.100 ;
        RECT 119.800 170.800 120.200 173.100 ;
        RECT 121.400 170.800 121.800 173.100 ;
        RECT 122.200 170.800 122.600 172.100 ;
        RECT 123.800 170.800 124.200 172.100 ;
        RECT 125.400 170.800 125.800 172.100 ;
        RECT 126.200 170.800 126.600 172.100 ;
        RECT 127.800 170.800 128.200 172.100 ;
        RECT 129.400 170.800 129.800 173.100 ;
        RECT 130.200 170.800 130.600 172.100 ;
        RECT 133.400 170.800 133.800 173.100 ;
        RECT 139.000 170.800 139.400 172.100 ;
        RECT 140.600 170.800 141.000 172.100 ;
        RECT 145.400 170.800 145.800 173.100 ;
        RECT 151.000 170.800 151.400 173.100 ;
        RECT 155.800 170.800 156.200 172.100 ;
        RECT 157.400 170.800 157.800 172.100 ;
        RECT 163.000 170.800 163.400 173.100 ;
        RECT 166.200 170.800 166.600 172.100 ;
        RECT 167.000 170.800 167.400 173.100 ;
        RECT 168.600 170.800 169.000 173.100 ;
        RECT 170.200 170.800 170.600 173.100 ;
        RECT 171.800 170.800 172.200 173.100 ;
        RECT 173.400 170.800 173.800 173.100 ;
        RECT 175.800 170.800 176.200 173.100 ;
        RECT 180.600 170.800 181.000 172.100 ;
        RECT 182.200 170.800 182.600 172.100 ;
        RECT 187.800 170.800 188.200 173.100 ;
        RECT 191.000 170.800 191.400 172.100 ;
        RECT 192.600 170.800 193.000 172.100 ;
        RECT 193.400 170.800 193.800 174.100 ;
        RECT 196.600 170.800 197.000 172.100 ;
        RECT 199.000 170.800 199.400 173.100 ;
        RECT 200.600 170.800 201.000 172.100 ;
        RECT 203.000 170.800 203.400 173.100 ;
        RECT 0.200 170.200 205.400 170.800 ;
        RECT 0.600 168.900 1.000 170.200 ;
        RECT 3.800 167.900 4.200 170.200 ;
        RECT 9.400 168.900 9.800 170.200 ;
        RECT 11.000 168.900 11.400 170.200 ;
        RECT 15.800 167.900 16.200 170.200 ;
        RECT 18.200 168.900 18.600 170.200 ;
        RECT 21.400 167.900 21.800 170.200 ;
        RECT 27.000 168.900 27.400 170.200 ;
        RECT 28.600 168.900 29.000 170.200 ;
        RECT 33.400 167.900 33.800 170.200 ;
        RECT 35.800 168.900 36.200 170.200 ;
        RECT 39.000 167.900 39.400 170.200 ;
        RECT 44.600 168.900 45.000 170.200 ;
        RECT 46.200 168.900 46.600 170.200 ;
        RECT 51.000 167.900 51.400 170.200 ;
        RECT 55.000 167.900 55.400 170.200 ;
        RECT 56.600 167.900 57.000 170.200 ;
        RECT 59.000 168.300 59.400 170.200 ;
        RECT 63.000 167.900 63.400 170.200 ;
        RECT 64.100 167.900 64.500 170.200 ;
        RECT 66.200 168.900 66.600 170.200 ;
        RECT 67.000 168.900 67.400 170.200 ;
        RECT 68.600 168.900 69.000 170.200 ;
        RECT 70.200 167.900 70.600 170.200 ;
        RECT 72.900 168.900 73.400 170.200 ;
        RECT 74.600 168.900 75.000 170.200 ;
        RECT 77.400 168.000 77.800 170.200 ;
        RECT 79.800 168.300 80.200 170.200 ;
        RECT 83.800 167.900 84.200 170.200 ;
        RECT 85.400 168.000 85.800 170.200 ;
        RECT 88.200 168.900 88.600 170.200 ;
        RECT 89.800 168.900 90.300 170.200 ;
        RECT 92.600 167.900 93.000 170.200 ;
        RECT 95.100 169.900 95.500 170.200 ;
        RECT 95.000 168.200 95.500 169.900 ;
        RECT 98.100 168.200 98.600 170.200 ;
        RECT 100.600 167.900 101.000 170.200 ;
        RECT 103.000 168.900 103.400 170.200 ;
        RECT 104.600 168.900 105.000 170.200 ;
        RECT 105.400 167.900 105.800 170.200 ;
        RECT 107.800 168.900 108.200 170.200 ;
        RECT 109.400 168.900 109.800 170.200 ;
        RECT 110.200 168.900 110.600 170.200 ;
        RECT 111.800 168.900 112.200 170.200 ;
        RECT 114.200 167.900 114.600 170.200 ;
        RECT 115.000 166.900 115.400 170.200 ;
        RECT 119.000 168.300 119.400 170.200 ;
        RECT 121.400 168.900 121.800 170.200 ;
        RECT 123.000 168.900 123.400 170.200 ;
        RECT 123.800 168.900 124.200 170.200 ;
        RECT 125.400 168.900 125.800 170.200 ;
        RECT 127.800 168.300 128.200 170.200 ;
        RECT 130.300 169.900 130.700 170.200 ;
        RECT 130.200 168.200 130.700 169.900 ;
        RECT 133.300 168.200 133.800 170.200 ;
        RECT 135.000 168.900 135.400 170.200 ;
        RECT 138.200 167.900 138.600 170.200 ;
        RECT 143.800 168.900 144.200 170.200 ;
        RECT 145.400 168.900 145.800 170.200 ;
        RECT 150.200 167.900 150.600 170.200 ;
        RECT 155.000 168.200 155.500 170.200 ;
        RECT 158.100 169.900 158.500 170.200 ;
        RECT 160.700 169.900 161.100 170.200 ;
        RECT 158.100 168.200 158.600 169.900 ;
        RECT 160.600 168.200 161.100 169.900 ;
        RECT 163.700 168.200 164.200 170.200 ;
        RECT 167.000 167.900 167.400 170.200 ;
        RECT 171.800 168.900 172.200 170.200 ;
        RECT 173.400 168.900 173.800 170.200 ;
        RECT 179.000 167.900 179.400 170.200 ;
        RECT 182.200 168.900 182.600 170.200 ;
        RECT 183.000 167.900 183.400 170.200 ;
        RECT 187.000 168.300 187.400 170.200 ;
        RECT 188.900 167.900 189.300 170.200 ;
        RECT 191.000 168.900 191.400 170.200 ;
        RECT 192.700 169.900 193.100 170.200 ;
        RECT 192.600 168.200 193.100 169.900 ;
        RECT 195.700 168.200 196.200 170.200 ;
        RECT 198.200 168.300 198.600 170.200 ;
        RECT 200.600 166.900 201.000 170.200 ;
        RECT 204.600 168.900 205.000 170.200 ;
        RECT 1.400 150.800 1.800 153.100 ;
        RECT 3.800 150.800 4.200 153.100 ;
        RECT 6.200 150.800 6.600 153.100 ;
        RECT 8.900 150.800 9.400 152.100 ;
        RECT 10.600 150.800 11.000 152.100 ;
        RECT 13.400 150.800 13.800 153.000 ;
        RECT 15.000 150.800 15.400 152.100 ;
        RECT 16.600 150.800 17.000 152.100 ;
        RECT 17.400 150.800 17.800 152.100 ;
        RECT 20.600 150.800 21.000 153.100 ;
        RECT 26.200 150.800 26.600 152.100 ;
        RECT 27.800 150.800 28.200 152.100 ;
        RECT 32.600 150.800 33.000 153.100 ;
        RECT 35.300 150.800 35.700 153.100 ;
        RECT 37.400 150.800 37.800 152.100 ;
        RECT 38.200 150.800 38.600 152.100 ;
        RECT 39.800 150.800 40.200 152.100 ;
        RECT 41.400 150.800 41.800 153.100 ;
        RECT 44.100 150.800 44.600 152.100 ;
        RECT 45.800 150.800 46.200 152.100 ;
        RECT 48.600 150.800 49.000 153.000 ;
        RECT 52.600 150.800 53.000 152.700 ;
        RECT 55.000 150.800 55.400 153.100 ;
        RECT 57.700 150.800 58.100 153.100 ;
        RECT 59.800 150.800 60.200 152.100 ;
        RECT 61.400 150.800 61.800 153.100 ;
        RECT 64.100 150.800 64.600 152.100 ;
        RECT 65.800 150.800 66.200 152.100 ;
        RECT 68.600 150.800 69.000 153.000 ;
        RECT 71.000 150.800 71.400 152.700 ;
        RECT 75.000 150.800 75.400 153.100 ;
        RECT 75.800 150.800 76.200 153.100 ;
        RECT 79.800 150.800 80.200 153.100 ;
        RECT 84.600 150.800 85.000 152.100 ;
        RECT 86.200 150.800 86.600 152.100 ;
        RECT 91.800 150.800 92.200 153.100 ;
        RECT 95.000 150.800 95.400 152.100 ;
        RECT 97.400 150.800 97.800 152.700 ;
        RECT 99.000 150.800 99.400 152.100 ;
        RECT 100.600 150.800 101.000 152.100 ;
        RECT 103.000 150.800 103.400 152.100 ;
        RECT 104.600 150.800 105.000 152.100 ;
        RECT 106.200 150.800 106.600 152.100 ;
        RECT 107.000 150.800 107.400 153.100 ;
        RECT 109.400 150.800 109.800 152.100 ;
        RECT 111.000 150.800 111.400 152.100 ;
        RECT 112.600 150.800 113.000 153.100 ;
        RECT 114.200 150.800 114.600 153.100 ;
        RECT 115.000 150.800 115.400 153.100 ;
        RECT 117.400 150.800 117.800 152.100 ;
        RECT 119.000 150.800 119.400 152.100 ;
        RECT 119.800 150.800 120.200 153.100 ;
        RECT 122.200 150.800 122.600 153.100 ;
        RECT 124.600 150.800 125.000 152.100 ;
        RECT 127.800 150.800 128.200 153.100 ;
        RECT 133.400 150.800 133.800 152.100 ;
        RECT 135.000 150.800 135.400 152.100 ;
        RECT 139.800 150.800 140.200 153.100 ;
        RECT 142.200 150.800 142.600 152.100 ;
        RECT 145.400 150.800 145.800 153.100 ;
        RECT 151.000 150.800 151.400 152.100 ;
        RECT 152.600 150.800 153.000 152.100 ;
        RECT 157.400 150.800 157.800 153.100 ;
        RECT 163.000 150.800 163.400 153.100 ;
        RECT 167.800 150.800 168.200 152.100 ;
        RECT 169.400 150.800 169.800 152.100 ;
        RECT 175.000 150.800 175.400 153.100 ;
        RECT 178.200 150.800 178.600 152.100 ;
        RECT 179.000 150.800 179.400 152.100 ;
        RECT 180.600 150.800 181.000 152.100 ;
        RECT 181.400 150.800 181.800 152.100 ;
        RECT 183.000 150.800 183.400 152.100 ;
        RECT 184.600 150.800 185.000 152.700 ;
        RECT 187.000 150.800 187.400 152.100 ;
        RECT 189.400 150.800 189.800 152.700 ;
        RECT 192.900 150.800 193.300 153.000 ;
        RECT 195.800 150.800 196.200 153.100 ;
        RECT 198.500 150.800 199.000 152.100 ;
        RECT 200.200 150.800 200.600 152.100 ;
        RECT 203.000 150.800 203.400 153.000 ;
        RECT 0.200 150.200 205.400 150.800 ;
        RECT 1.400 147.900 1.800 150.200 ;
        RECT 4.100 148.900 4.600 150.200 ;
        RECT 5.800 148.900 6.200 150.200 ;
        RECT 8.600 148.000 9.000 150.200 ;
        RECT 11.000 148.300 11.400 150.200 ;
        RECT 13.700 147.900 14.100 150.200 ;
        RECT 15.800 148.900 16.200 150.200 ;
        RECT 16.600 147.900 17.000 150.200 ;
        RECT 20.600 148.300 21.000 150.200 ;
        RECT 23.000 147.900 23.400 150.200 ;
        RECT 25.700 148.900 26.200 150.200 ;
        RECT 27.400 148.900 27.800 150.200 ;
        RECT 30.200 148.000 30.600 150.200 ;
        RECT 32.600 147.900 33.000 150.200 ;
        RECT 35.300 148.900 35.800 150.200 ;
        RECT 37.000 148.900 37.400 150.200 ;
        RECT 39.800 148.000 40.200 150.200 ;
        RECT 42.200 147.900 42.600 150.200 ;
        RECT 44.900 148.900 45.400 150.200 ;
        RECT 46.600 148.900 47.000 150.200 ;
        RECT 49.400 148.000 49.800 150.200 ;
        RECT 53.400 148.900 53.800 150.200 ;
        RECT 54.200 147.900 54.600 150.200 ;
        RECT 58.200 148.300 58.600 150.200 ;
        RECT 60.600 147.900 61.000 150.200 ;
        RECT 62.200 147.900 62.600 150.200 ;
        RECT 63.000 148.900 63.400 150.200 ;
        RECT 64.600 148.900 65.000 150.200 ;
        RECT 66.200 148.900 66.600 150.200 ;
        RECT 67.000 148.900 67.400 150.200 ;
        RECT 70.200 147.900 70.600 150.200 ;
        RECT 75.800 148.900 76.200 150.200 ;
        RECT 77.400 148.900 77.800 150.200 ;
        RECT 82.200 147.900 82.600 150.200 ;
        RECT 84.600 148.900 85.000 150.200 ;
        RECT 87.000 148.300 87.400 150.200 ;
        RECT 91.000 147.900 91.400 150.200 ;
        RECT 92.600 148.000 93.000 150.200 ;
        RECT 95.400 148.900 95.800 150.200 ;
        RECT 97.000 148.900 97.500 150.200 ;
        RECT 99.800 147.900 100.200 150.200 ;
        RECT 105.400 146.900 105.800 150.200 ;
        RECT 106.200 146.900 106.600 150.200 ;
        RECT 109.400 148.900 109.800 150.200 ;
        RECT 111.000 148.900 111.400 150.200 ;
        RECT 113.400 147.900 113.800 150.200 ;
        RECT 114.200 146.900 114.600 150.200 ;
        RECT 117.400 146.900 117.800 150.200 ;
        RECT 120.600 146.900 121.000 150.200 ;
        RECT 123.800 146.900 124.200 150.200 ;
        RECT 127.000 146.900 127.400 150.200 ;
        RECT 130.200 148.900 130.600 150.200 ;
        RECT 131.800 148.900 132.200 150.200 ;
        RECT 132.600 147.900 133.000 150.200 ;
        RECT 134.200 147.900 134.600 150.200 ;
        RECT 135.800 148.900 136.200 150.200 ;
        RECT 137.400 148.900 137.800 150.200 ;
        RECT 139.000 148.200 139.500 150.200 ;
        RECT 142.100 149.900 142.500 150.200 ;
        RECT 142.100 148.200 142.600 149.900 ;
        RECT 143.800 147.900 144.200 150.200 ;
        RECT 146.200 147.900 146.600 150.200 ;
        RECT 148.900 147.900 149.300 150.200 ;
        RECT 151.000 148.900 151.400 150.200 ;
        RECT 153.400 147.900 153.800 150.200 ;
        RECT 156.400 147.900 156.800 150.200 ;
        RECT 159.000 148.300 159.400 150.200 ;
        RECT 160.600 148.900 161.000 150.200 ;
        RECT 162.200 147.900 162.600 150.200 ;
        RECT 165.400 148.300 165.800 150.200 ;
        RECT 167.800 147.900 168.200 150.200 ;
        RECT 170.800 147.900 171.200 150.200 ;
        RECT 171.800 147.900 172.200 150.200 ;
        RECT 174.200 148.900 174.600 150.200 ;
        RECT 176.300 147.900 176.700 150.200 ;
        RECT 177.400 147.900 177.800 150.200 ;
        RECT 179.800 148.900 180.200 150.200 ;
        RECT 181.400 148.900 181.800 150.200 ;
        RECT 182.400 147.900 182.800 150.200 ;
        RECT 185.400 147.900 185.800 150.200 ;
        RECT 186.200 148.900 186.600 150.200 ;
        RECT 187.800 148.900 188.200 150.200 ;
        RECT 188.600 147.900 189.000 150.200 ;
        RECT 191.000 148.900 191.400 150.200 ;
        RECT 192.600 148.900 193.000 150.200 ;
        RECT 193.400 146.900 193.800 150.200 ;
        RECT 199.000 146.900 199.400 150.200 ;
        RECT 200.900 148.000 201.300 150.200 ;
        RECT 203.800 147.900 204.200 150.200 ;
        RECT 0.600 130.800 1.000 132.100 ;
        RECT 3.800 130.800 4.200 133.100 ;
        RECT 9.400 130.800 9.800 132.100 ;
        RECT 11.000 130.800 11.400 132.100 ;
        RECT 15.800 130.800 16.200 133.100 ;
        RECT 19.800 130.800 20.200 133.100 ;
        RECT 20.600 130.800 21.000 132.100 ;
        RECT 23.800 130.800 24.200 133.100 ;
        RECT 29.400 130.800 29.800 132.100 ;
        RECT 31.000 130.800 31.400 132.100 ;
        RECT 35.800 130.800 36.200 133.100 ;
        RECT 39.000 130.800 39.400 132.700 ;
        RECT 41.700 130.800 42.100 133.100 ;
        RECT 43.800 130.800 44.200 132.100 ;
        RECT 46.200 130.800 46.600 132.700 ;
        RECT 47.800 130.800 48.200 132.100 ;
        RECT 49.900 130.800 50.300 133.100 ;
        RECT 53.400 130.800 53.800 133.100 ;
        RECT 56.100 130.800 56.600 132.100 ;
        RECT 57.800 130.800 58.200 132.100 ;
        RECT 60.600 130.800 61.000 133.000 ;
        RECT 62.200 130.800 62.600 133.100 ;
        RECT 66.200 130.800 66.600 132.700 ;
        RECT 68.600 130.800 69.000 132.700 ;
        RECT 72.600 130.800 73.000 133.100 ;
        RECT 73.700 130.800 74.100 133.100 ;
        RECT 75.800 130.800 76.200 132.100 ;
        RECT 76.600 130.800 77.000 133.100 ;
        RECT 80.600 130.800 81.000 132.700 ;
        RECT 83.000 130.800 83.400 133.000 ;
        RECT 85.800 130.800 86.200 132.100 ;
        RECT 87.400 130.800 87.900 132.100 ;
        RECT 90.200 130.800 90.600 133.100 ;
        RECT 91.800 130.800 92.200 133.100 ;
        RECT 95.800 130.800 96.200 132.700 ;
        RECT 97.400 130.800 97.800 133.100 ;
        RECT 99.000 130.800 99.400 133.100 ;
        RECT 103.000 130.800 103.400 133.100 ;
        RECT 104.600 130.800 105.000 133.100 ;
        RECT 106.200 130.800 106.600 133.300 ;
        RECT 108.800 130.800 109.200 133.500 ;
        RECT 111.000 130.800 111.400 132.700 ;
        RECT 115.000 130.800 115.400 133.100 ;
        RECT 116.600 130.800 117.000 133.000 ;
        RECT 119.400 130.800 119.800 132.100 ;
        RECT 121.000 130.800 121.500 132.100 ;
        RECT 123.800 130.800 124.200 133.100 ;
        RECT 127.000 130.800 127.400 133.100 ;
        RECT 127.800 130.800 128.200 133.100 ;
        RECT 130.200 130.800 130.600 132.100 ;
        RECT 131.800 130.800 132.200 132.100 ;
        RECT 132.600 130.800 133.000 132.100 ;
        RECT 134.200 130.800 134.600 132.100 ;
        RECT 135.000 130.800 135.400 132.100 ;
        RECT 136.600 130.800 137.000 132.100 ;
        RECT 137.400 130.800 137.800 132.100 ;
        RECT 139.500 130.800 139.900 133.100 ;
        RECT 140.600 130.800 141.000 133.100 ;
        RECT 142.200 130.800 142.600 133.100 ;
        RECT 144.600 130.800 145.000 133.100 ;
        RECT 146.200 130.800 146.600 133.100 ;
        RECT 147.800 130.800 148.200 133.100 ;
        RECT 149.400 130.800 149.800 133.100 ;
        RECT 152.600 130.800 153.000 133.100 ;
        RECT 155.300 130.800 155.800 132.100 ;
        RECT 157.000 130.800 157.400 132.100 ;
        RECT 159.800 130.800 160.200 133.000 ;
        RECT 161.400 130.800 161.800 132.100 ;
        RECT 163.000 130.800 163.400 132.100 ;
        RECT 163.800 130.800 164.200 132.100 ;
        RECT 166.200 130.800 166.600 133.300 ;
        RECT 168.800 130.800 169.200 133.500 ;
        RECT 171.800 130.800 172.200 133.100 ;
        RECT 174.200 130.800 174.600 132.700 ;
        RECT 178.200 130.800 178.600 134.100 ;
        RECT 179.000 130.800 179.400 133.100 ;
        RECT 182.500 130.800 182.900 133.000 ;
        RECT 186.200 130.800 186.600 132.700 ;
        RECT 189.400 130.800 189.800 133.100 ;
        RECT 191.800 130.800 192.200 133.100 ;
        RECT 195.000 130.800 195.400 134.100 ;
        RECT 195.800 130.800 196.200 132.100 ;
        RECT 197.900 130.800 198.300 133.100 ;
        RECT 199.800 130.800 200.300 132.800 ;
        RECT 202.900 131.100 203.400 132.800 ;
        RECT 202.900 130.800 203.300 131.100 ;
        RECT 0.200 130.200 205.400 130.800 ;
        RECT 1.400 127.900 1.800 130.200 ;
        RECT 4.100 128.900 4.600 130.200 ;
        RECT 5.800 128.900 6.200 130.200 ;
        RECT 8.600 128.000 9.000 130.200 ;
        RECT 10.200 128.900 10.600 130.200 ;
        RECT 12.400 127.500 12.800 130.200 ;
        RECT 15.000 127.700 15.400 130.200 ;
        RECT 17.400 127.900 17.800 130.200 ;
        RECT 20.100 128.900 20.600 130.200 ;
        RECT 21.800 128.900 22.200 130.200 ;
        RECT 24.600 128.000 25.000 130.200 ;
        RECT 27.000 128.300 27.400 130.200 ;
        RECT 31.000 127.900 31.400 130.200 ;
        RECT 32.600 127.900 33.000 130.200 ;
        RECT 35.300 128.900 35.800 130.200 ;
        RECT 37.000 128.900 37.400 130.200 ;
        RECT 39.800 128.000 40.200 130.200 ;
        RECT 41.400 127.900 41.800 130.200 ;
        RECT 44.600 128.300 45.000 130.200 ;
        RECT 47.800 128.300 48.200 130.200 ;
        RECT 52.900 127.900 53.300 130.200 ;
        RECT 55.000 128.900 55.400 130.200 ;
        RECT 57.400 128.300 57.800 130.200 ;
        RECT 60.600 127.900 61.000 130.200 ;
        RECT 61.400 128.900 61.800 130.200 ;
        RECT 64.600 128.300 65.000 130.200 ;
        RECT 67.000 128.300 67.400 130.200 ;
        RECT 70.200 128.300 70.600 130.200 ;
        RECT 73.400 128.000 73.800 130.200 ;
        RECT 76.200 128.900 76.600 130.200 ;
        RECT 77.800 128.900 78.300 130.200 ;
        RECT 80.600 127.900 81.000 130.200 ;
        RECT 83.800 128.300 84.200 130.200 ;
        RECT 85.400 128.900 85.800 130.200 ;
        RECT 87.000 128.900 87.400 130.200 ;
        RECT 88.600 128.900 89.000 130.200 ;
        RECT 90.200 128.000 90.600 130.200 ;
        RECT 93.000 128.900 93.400 130.200 ;
        RECT 94.600 128.900 95.100 130.200 ;
        RECT 97.400 127.900 97.800 130.200 ;
        RECT 99.000 127.900 99.400 130.200 ;
        RECT 104.600 128.300 105.000 130.200 ;
        RECT 107.800 128.300 108.200 130.200 ;
        RECT 111.800 128.300 112.200 130.200 ;
        RECT 113.400 128.900 113.800 130.200 ;
        RECT 115.000 128.900 115.400 130.200 ;
        RECT 115.800 128.900 116.200 130.200 ;
        RECT 117.400 128.900 117.800 130.200 ;
        RECT 119.000 128.000 119.400 130.200 ;
        RECT 121.800 128.900 122.200 130.200 ;
        RECT 123.400 128.900 123.900 130.200 ;
        RECT 126.200 127.900 126.600 130.200 ;
        RECT 128.600 127.900 129.000 130.200 ;
        RECT 131.300 128.900 131.800 130.200 ;
        RECT 133.000 128.900 133.400 130.200 ;
        RECT 135.800 128.000 136.200 130.200 ;
        RECT 138.200 128.300 138.600 130.200 ;
        RECT 142.200 127.900 142.600 130.200 ;
        RECT 143.000 128.900 143.400 130.200 ;
        RECT 145.400 128.000 145.800 130.200 ;
        RECT 148.200 128.900 148.600 130.200 ;
        RECT 149.800 128.900 150.300 130.200 ;
        RECT 152.600 127.900 153.000 130.200 ;
        RECT 155.800 128.900 156.200 130.200 ;
        RECT 157.400 128.900 157.800 130.200 ;
        RECT 158.200 128.900 158.600 130.200 ;
        RECT 160.300 127.900 160.700 130.200 ;
        RECT 161.400 128.900 161.800 130.200 ;
        RECT 163.500 127.900 163.900 130.200 ;
        RECT 166.200 128.300 166.600 130.200 ;
        RECT 168.100 127.900 168.500 130.200 ;
        RECT 170.200 128.900 170.600 130.200 ;
        RECT 172.600 128.300 173.000 130.200 ;
        RECT 175.000 127.900 175.400 130.200 ;
        RECT 176.600 127.900 177.000 130.200 ;
        RECT 179.000 127.900 179.400 130.200 ;
        RECT 181.400 127.900 181.800 130.200 ;
        RECT 183.000 127.900 183.400 130.200 ;
        RECT 184.600 127.900 185.000 130.200 ;
        RECT 185.400 127.900 185.800 130.200 ;
        RECT 187.000 127.900 187.400 130.200 ;
        RECT 187.800 127.900 188.200 130.200 ;
        RECT 189.400 127.900 189.800 130.200 ;
        RECT 190.200 127.900 190.600 130.200 ;
        RECT 191.800 127.900 192.200 130.200 ;
        RECT 193.400 127.700 193.800 130.200 ;
        RECT 196.000 127.500 196.400 130.200 ;
        RECT 197.700 127.900 198.100 130.200 ;
        RECT 199.800 128.900 200.200 130.200 ;
        RECT 201.400 128.900 201.800 130.200 ;
        RECT 202.200 128.900 202.600 130.200 ;
        RECT 203.800 128.900 204.200 130.200 ;
        RECT 1.400 110.800 1.800 113.100 ;
        RECT 4.100 110.800 4.600 112.100 ;
        RECT 5.800 110.800 6.200 112.100 ;
        RECT 8.600 110.800 9.000 113.000 ;
        RECT 11.000 110.800 11.400 113.100 ;
        RECT 13.700 110.800 14.200 112.100 ;
        RECT 15.400 110.800 15.800 112.100 ;
        RECT 18.200 110.800 18.600 113.000 ;
        RECT 19.800 110.800 20.200 112.100 ;
        RECT 22.200 110.800 22.600 113.300 ;
        RECT 24.800 110.800 25.200 113.500 ;
        RECT 27.000 110.800 27.400 113.100 ;
        RECT 29.700 110.800 30.200 112.100 ;
        RECT 31.400 110.800 31.800 112.100 ;
        RECT 34.200 110.800 34.600 113.000 ;
        RECT 35.800 110.800 36.200 113.100 ;
        RECT 39.800 110.800 40.200 112.700 ;
        RECT 42.200 110.800 42.600 112.700 ;
        RECT 44.600 110.800 45.000 112.100 ;
        RECT 46.700 110.800 47.100 113.100 ;
        RECT 47.800 110.800 48.200 113.100 ;
        RECT 49.400 110.800 49.800 113.100 ;
        RECT 53.400 110.800 53.800 112.700 ;
        RECT 57.400 110.800 57.800 113.100 ;
        RECT 58.200 110.800 58.600 112.100 ;
        RECT 60.300 110.800 60.700 113.100 ;
        RECT 62.200 110.800 62.600 112.700 ;
        RECT 65.400 110.800 65.800 113.000 ;
        RECT 68.200 110.800 68.600 112.100 ;
        RECT 69.800 110.800 70.300 112.100 ;
        RECT 72.600 110.800 73.000 113.100 ;
        RECT 74.200 110.800 74.600 113.100 ;
        RECT 75.800 110.800 76.200 113.100 ;
        RECT 78.200 110.800 78.600 113.100 ;
        RECT 79.800 110.800 80.200 113.100 ;
        RECT 81.400 110.800 81.800 113.100 ;
        RECT 83.000 110.800 83.400 113.100 ;
        RECT 83.800 110.800 84.200 112.100 ;
        RECT 85.900 110.800 86.300 113.100 ;
        RECT 87.800 110.800 88.200 112.700 ;
        RECT 90.200 110.800 90.600 113.100 ;
        RECT 93.400 110.800 93.800 113.100 ;
        RECT 96.100 110.800 96.600 112.100 ;
        RECT 97.800 110.800 98.200 112.100 ;
        RECT 100.600 110.800 101.000 113.000 ;
        RECT 103.800 110.800 104.200 113.100 ;
        RECT 107.800 110.800 108.200 112.700 ;
        RECT 110.200 110.800 110.600 113.100 ;
        RECT 111.800 110.800 112.200 113.100 ;
        RECT 113.400 110.800 113.900 112.800 ;
        RECT 116.500 111.100 117.000 112.800 ;
        RECT 116.500 110.800 116.900 111.100 ;
        RECT 118.200 110.800 118.600 113.100 ;
        RECT 119.800 110.800 120.200 113.100 ;
        RECT 123.000 110.800 123.400 112.700 ;
        RECT 124.900 110.800 125.300 113.100 ;
        RECT 127.000 110.800 127.400 112.100 ;
        RECT 129.400 110.800 129.800 112.700 ;
        RECT 131.000 110.800 131.400 113.100 ;
        RECT 133.400 110.800 133.800 112.100 ;
        RECT 136.600 110.800 137.000 113.100 ;
        RECT 142.200 110.800 142.600 112.100 ;
        RECT 143.800 110.800 144.200 112.100 ;
        RECT 148.600 110.800 149.000 113.100 ;
        RECT 151.000 110.800 151.400 112.100 ;
        RECT 152.600 110.800 153.000 112.100 ;
        RECT 155.000 110.800 155.400 112.100 ;
        RECT 157.100 110.800 157.500 113.100 ;
        RECT 158.200 110.800 158.600 112.100 ;
        RECT 160.300 110.800 160.700 113.100 ;
        RECT 163.800 110.800 164.200 114.100 ;
        RECT 165.400 110.800 165.800 112.700 ;
        RECT 169.400 110.800 169.800 113.100 ;
        RECT 174.200 110.800 174.600 112.100 ;
        RECT 175.800 110.800 176.200 112.100 ;
        RECT 181.400 110.800 181.800 113.100 ;
        RECT 184.600 110.800 185.000 112.100 ;
        RECT 186.200 110.800 186.600 113.000 ;
        RECT 189.000 110.800 189.400 112.100 ;
        RECT 190.600 110.800 191.100 112.100 ;
        RECT 193.400 110.800 193.800 113.100 ;
        RECT 195.800 110.800 196.200 113.100 ;
        RECT 198.500 110.800 199.000 112.100 ;
        RECT 200.200 110.800 200.600 112.100 ;
        RECT 203.000 110.800 203.400 113.000 ;
        RECT 0.200 110.200 205.400 110.800 ;
        RECT 1.400 108.000 1.800 110.200 ;
        RECT 4.200 108.900 4.600 110.200 ;
        RECT 5.800 108.900 6.300 110.200 ;
        RECT 8.600 107.900 9.000 110.200 ;
        RECT 10.200 108.900 10.600 110.200 ;
        RECT 12.600 108.300 13.000 110.200 ;
        RECT 16.600 107.900 17.000 110.200 ;
        RECT 18.000 107.500 18.400 110.200 ;
        RECT 20.600 107.700 21.000 110.200 ;
        RECT 22.200 108.900 22.600 110.200 ;
        RECT 24.600 108.300 25.000 110.200 ;
        RECT 27.000 108.900 27.400 110.200 ;
        RECT 28.900 107.900 29.300 110.200 ;
        RECT 31.000 108.900 31.400 110.200 ;
        RECT 33.400 108.300 33.800 110.200 ;
        RECT 35.000 108.900 35.400 110.200 ;
        RECT 37.400 108.300 37.800 110.200 ;
        RECT 39.800 108.900 40.200 110.200 ;
        RECT 41.900 107.900 42.300 110.200 ;
        RECT 43.300 107.900 43.700 110.200 ;
        RECT 45.400 108.900 45.800 110.200 ;
        RECT 46.200 107.900 46.600 110.200 ;
        RECT 47.800 107.900 48.200 110.200 ;
        RECT 51.800 107.900 52.200 110.200 ;
        RECT 53.400 107.900 53.800 110.200 ;
        RECT 54.200 107.900 54.600 110.200 ;
        RECT 55.800 107.900 56.200 110.200 ;
        RECT 59.800 108.300 60.200 110.200 ;
        RECT 61.400 107.900 61.800 110.200 ;
        RECT 63.000 107.900 63.400 110.200 ;
        RECT 64.600 108.900 65.000 110.200 ;
        RECT 66.200 108.900 66.600 110.200 ;
        RECT 68.300 107.900 68.700 110.200 ;
        RECT 70.200 108.300 70.600 110.200 ;
        RECT 73.400 108.900 73.800 110.200 ;
        RECT 75.000 108.900 75.400 110.200 ;
        RECT 76.600 107.900 77.000 110.200 ;
        RECT 79.300 108.900 79.800 110.200 ;
        RECT 81.000 108.900 81.400 110.200 ;
        RECT 83.800 108.000 84.200 110.200 ;
        RECT 87.000 107.900 87.400 110.200 ;
        RECT 87.800 108.900 88.200 110.200 ;
        RECT 89.400 108.900 89.800 110.200 ;
        RECT 91.800 108.300 92.200 110.200 ;
        RECT 93.400 107.900 93.800 110.200 ;
        RECT 95.000 107.900 95.400 110.200 ;
        RECT 97.400 108.900 97.800 110.200 ;
        RECT 98.200 107.900 98.600 110.200 ;
        RECT 103.800 108.300 104.200 110.200 ;
        RECT 106.200 108.000 106.600 110.200 ;
        RECT 109.000 108.900 109.400 110.200 ;
        RECT 110.600 108.900 111.100 110.200 ;
        RECT 113.400 107.900 113.800 110.200 ;
        RECT 115.800 107.900 116.200 110.200 ;
        RECT 117.400 107.900 117.800 110.200 ;
        RECT 119.000 107.900 119.400 110.200 ;
        RECT 121.700 108.900 122.200 110.200 ;
        RECT 123.400 108.900 123.800 110.200 ;
        RECT 126.200 108.000 126.600 110.200 ;
        RECT 127.800 108.900 128.200 110.200 ;
        RECT 129.400 108.900 129.800 110.200 ;
        RECT 130.200 108.900 130.600 110.200 ;
        RECT 132.300 107.900 132.700 110.200 ;
        RECT 134.200 107.700 134.600 110.200 ;
        RECT 136.800 107.500 137.200 110.200 ;
        RECT 139.000 108.900 139.400 110.200 ;
        RECT 140.600 108.000 141.000 110.200 ;
        RECT 143.400 108.900 143.800 110.200 ;
        RECT 145.000 108.900 145.500 110.200 ;
        RECT 147.800 107.900 148.200 110.200 ;
        RECT 151.800 107.900 152.200 110.200 ;
        RECT 154.500 108.900 155.000 110.200 ;
        RECT 156.200 108.900 156.600 110.200 ;
        RECT 159.000 108.000 159.400 110.200 ;
        RECT 160.900 107.900 161.300 110.200 ;
        RECT 163.000 108.900 163.400 110.200 ;
        RECT 163.800 108.900 164.200 110.200 ;
        RECT 165.400 108.900 165.800 110.200 ;
        RECT 166.500 107.900 166.900 110.200 ;
        RECT 168.600 108.900 169.000 110.200 ;
        RECT 170.200 107.900 170.600 110.200 ;
        RECT 171.800 107.900 172.200 110.200 ;
        RECT 174.200 108.300 174.600 110.200 ;
        RECT 176.600 108.900 177.000 110.200 ;
        RECT 178.200 108.000 178.600 110.200 ;
        RECT 181.000 108.900 181.400 110.200 ;
        RECT 182.600 108.900 183.100 110.200 ;
        RECT 185.400 107.900 185.800 110.200 ;
        RECT 187.800 107.700 188.200 110.200 ;
        RECT 190.400 107.500 190.800 110.200 ;
        RECT 192.600 107.700 193.000 110.200 ;
        RECT 195.200 107.500 195.600 110.200 ;
        RECT 197.400 108.300 197.800 110.200 ;
        RECT 201.400 107.900 201.800 110.200 ;
        RECT 203.800 107.900 204.200 110.200 ;
        RECT 0.600 90.800 1.000 93.100 ;
        RECT 2.200 90.800 2.600 93.100 ;
        RECT 3.800 90.800 4.200 93.100 ;
        RECT 5.400 90.800 5.800 93.100 ;
        RECT 7.000 90.800 7.400 93.100 ;
        RECT 8.600 90.800 9.000 93.100 ;
        RECT 11.300 90.800 11.800 92.100 ;
        RECT 13.000 90.800 13.400 92.100 ;
        RECT 15.800 90.800 16.200 93.000 ;
        RECT 18.200 90.800 18.600 92.700 ;
        RECT 20.600 90.800 21.000 93.100 ;
        RECT 23.300 90.800 23.700 93.100 ;
        RECT 25.400 90.800 25.800 92.100 ;
        RECT 26.200 90.800 26.600 92.100 ;
        RECT 28.100 90.800 28.500 93.100 ;
        RECT 30.200 90.800 30.600 92.100 ;
        RECT 31.300 90.800 31.700 93.100 ;
        RECT 33.400 90.800 33.800 92.100 ;
        RECT 35.000 90.800 35.400 92.700 ;
        RECT 38.200 90.800 38.600 92.700 ;
        RECT 40.600 90.800 41.000 92.100 ;
        RECT 42.700 90.800 43.100 93.100 ;
        RECT 45.400 90.800 45.800 92.700 ;
        RECT 47.800 90.800 48.200 92.700 ;
        RECT 52.600 90.800 53.000 93.100 ;
        RECT 54.200 90.800 54.600 93.100 ;
        RECT 57.400 90.800 57.800 92.700 ;
        RECT 59.300 90.800 59.700 93.100 ;
        RECT 61.400 90.800 61.800 92.100 ;
        RECT 62.200 90.800 62.600 92.100 ;
        RECT 64.300 90.800 64.700 93.100 ;
        RECT 66.200 90.800 66.600 93.100 ;
        RECT 67.800 90.800 68.200 93.100 ;
        RECT 68.600 90.800 69.000 93.100 ;
        RECT 70.200 90.800 70.600 93.100 ;
        RECT 71.800 90.800 72.200 93.100 ;
        RECT 75.000 90.800 75.400 92.700 ;
        RECT 78.200 90.800 78.600 92.700 ;
        RECT 81.400 90.800 81.800 92.700 ;
        RECT 84.600 90.800 85.000 92.700 ;
        RECT 87.000 90.800 87.400 92.700 ;
        RECT 90.200 90.800 90.600 92.100 ;
        RECT 92.300 90.800 92.700 93.100 ;
        RECT 95.000 90.800 95.400 92.700 ;
        RECT 96.600 90.800 97.000 93.100 ;
        RECT 98.200 90.800 98.600 93.100 ;
        RECT 99.800 90.800 100.200 93.100 ;
        RECT 101.400 90.800 101.800 93.100 ;
        RECT 105.400 90.800 105.800 93.100 ;
        RECT 108.100 90.800 108.600 92.100 ;
        RECT 109.800 90.800 110.200 92.100 ;
        RECT 112.600 90.800 113.000 93.000 ;
        RECT 115.000 90.800 115.400 92.700 ;
        RECT 117.400 90.800 117.800 93.100 ;
        RECT 121.400 90.800 121.800 92.700 ;
        RECT 123.000 90.800 123.400 93.100 ;
        RECT 124.600 90.800 125.000 93.100 ;
        RECT 127.000 90.800 127.400 93.100 ;
        RECT 128.600 90.800 129.000 93.100 ;
        RECT 130.200 90.800 130.600 93.100 ;
        RECT 132.900 90.800 133.400 92.100 ;
        RECT 134.600 90.800 135.000 92.100 ;
        RECT 137.400 90.800 137.800 93.000 ;
        RECT 139.300 90.800 139.700 93.100 ;
        RECT 141.400 90.800 141.800 92.100 ;
        RECT 142.200 90.800 142.600 92.100 ;
        RECT 143.800 90.800 144.200 92.100 ;
        RECT 145.400 90.800 145.800 92.700 ;
        RECT 148.100 90.800 148.500 93.100 ;
        RECT 150.200 90.800 150.600 92.100 ;
        RECT 151.800 90.800 152.200 93.100 ;
        RECT 153.400 90.800 153.800 93.100 ;
        RECT 156.600 90.800 157.000 92.900 ;
        RECT 158.200 90.800 158.600 92.100 ;
        RECT 159.000 90.800 159.400 92.100 ;
        RECT 161.100 90.800 161.500 93.100 ;
        RECT 162.200 90.800 162.600 93.100 ;
        RECT 166.200 90.800 166.600 92.700 ;
        RECT 169.400 90.800 169.800 92.700 ;
        RECT 171.800 90.800 172.200 92.700 ;
        RECT 174.200 90.800 174.600 92.100 ;
        RECT 176.300 90.800 176.700 93.100 ;
        RECT 178.200 90.800 178.600 93.300 ;
        RECT 180.800 90.800 181.200 93.500 ;
        RECT 183.000 90.800 183.400 92.100 ;
        RECT 184.600 90.800 185.000 93.000 ;
        RECT 187.400 90.800 187.800 92.100 ;
        RECT 189.000 90.800 189.500 92.100 ;
        RECT 191.800 90.800 192.200 93.100 ;
        RECT 194.200 90.800 194.600 92.100 ;
        RECT 195.800 90.800 196.200 93.000 ;
        RECT 198.600 90.800 199.000 92.100 ;
        RECT 200.200 90.800 200.700 92.100 ;
        RECT 203.000 90.800 203.400 93.100 ;
        RECT 0.200 90.200 205.400 90.800 ;
        RECT 1.400 88.000 1.800 90.200 ;
        RECT 4.200 88.900 4.600 90.200 ;
        RECT 5.800 88.900 6.300 90.200 ;
        RECT 8.600 87.900 9.000 90.200 ;
        RECT 10.200 87.900 10.600 90.200 ;
        RECT 14.200 88.300 14.600 90.200 ;
        RECT 17.400 87.900 17.800 90.200 ;
        RECT 18.500 87.900 18.900 90.200 ;
        RECT 20.600 88.900 21.000 90.200 ;
        RECT 23.000 88.300 23.400 90.200 ;
        RECT 25.400 87.900 25.800 90.200 ;
        RECT 28.100 88.900 28.600 90.200 ;
        RECT 29.800 88.900 30.200 90.200 ;
        RECT 32.600 88.000 33.000 90.200 ;
        RECT 34.200 88.900 34.600 90.200 ;
        RECT 35.800 88.900 36.200 90.200 ;
        RECT 36.600 88.900 37.000 90.200 ;
        RECT 38.700 87.900 39.100 90.200 ;
        RECT 40.100 87.900 40.500 90.200 ;
        RECT 42.200 88.900 42.600 90.200 ;
        RECT 44.600 88.300 45.000 90.200 ;
        RECT 47.000 88.900 47.400 90.200 ;
        RECT 50.200 88.000 50.600 90.200 ;
        RECT 53.000 88.900 53.400 90.200 ;
        RECT 54.600 88.900 55.100 90.200 ;
        RECT 57.400 87.900 57.800 90.200 ;
        RECT 59.000 87.900 59.400 90.200 ;
        RECT 63.000 88.300 63.400 90.200 ;
        RECT 65.400 87.900 65.800 90.200 ;
        RECT 67.000 87.900 67.400 90.200 ;
        RECT 69.400 88.300 69.800 90.200 ;
        RECT 72.600 88.300 73.000 90.200 ;
        RECT 74.200 88.900 74.600 90.200 ;
        RECT 76.300 87.900 76.700 90.200 ;
        RECT 77.400 87.900 77.800 90.200 ;
        RECT 79.000 87.900 79.400 90.200 ;
        RECT 81.400 88.300 81.800 90.200 ;
        RECT 85.400 88.300 85.800 90.200 ;
        RECT 87.000 87.900 87.400 90.200 ;
        RECT 88.600 87.900 89.000 90.200 ;
        RECT 90.200 87.900 90.600 90.200 ;
        RECT 91.300 87.900 91.700 90.200 ;
        RECT 93.400 88.900 93.800 90.200 ;
        RECT 95.800 88.300 96.200 90.200 ;
        RECT 98.200 88.900 98.600 90.200 ;
        RECT 99.000 87.900 99.400 90.200 ;
        RECT 104.600 88.300 105.000 90.200 ;
        RECT 107.000 88.000 107.400 90.200 ;
        RECT 109.800 88.900 110.200 90.200 ;
        RECT 111.400 88.900 111.900 90.200 ;
        RECT 114.200 87.900 114.600 90.200 ;
        RECT 115.800 88.900 116.200 90.200 ;
        RECT 117.900 87.900 118.300 90.200 ;
        RECT 119.800 88.000 120.200 90.200 ;
        RECT 122.600 88.900 123.000 90.200 ;
        RECT 124.200 88.900 124.700 90.200 ;
        RECT 127.000 87.900 127.400 90.200 ;
        RECT 128.600 88.900 129.000 90.200 ;
        RECT 130.200 88.900 130.600 90.200 ;
        RECT 131.000 88.900 131.400 90.200 ;
        RECT 133.100 87.900 133.500 90.200 ;
        RECT 135.000 87.900 135.400 90.200 ;
        RECT 136.600 87.900 137.000 90.200 ;
        RECT 138.200 88.000 138.600 90.200 ;
        RECT 141.000 88.900 141.400 90.200 ;
        RECT 142.600 88.900 143.100 90.200 ;
        RECT 145.400 87.900 145.800 90.200 ;
        RECT 148.600 88.300 149.000 90.200 ;
        RECT 151.000 87.700 151.400 90.200 ;
        RECT 153.600 87.500 154.000 90.200 ;
        RECT 156.600 88.900 157.000 90.200 ;
        RECT 158.700 87.900 159.100 90.200 ;
        RECT 160.600 88.900 161.000 90.200 ;
        RECT 162.200 88.000 162.600 90.200 ;
        RECT 165.000 88.900 165.400 90.200 ;
        RECT 166.600 88.900 167.100 90.200 ;
        RECT 169.400 87.900 169.800 90.200 ;
        RECT 171.800 88.300 172.200 90.200 ;
        RECT 175.800 87.900 176.200 90.200 ;
        RECT 178.200 88.300 178.600 90.200 ;
        RECT 180.600 88.000 181.000 90.200 ;
        RECT 183.400 88.900 183.800 90.200 ;
        RECT 185.000 88.900 185.500 90.200 ;
        RECT 187.800 87.900 188.200 90.200 ;
        RECT 190.000 87.500 190.400 90.200 ;
        RECT 192.600 87.700 193.000 90.200 ;
        RECT 195.000 88.900 195.400 90.200 ;
        RECT 196.600 88.000 197.000 90.200 ;
        RECT 199.400 88.900 199.800 90.200 ;
        RECT 201.000 88.900 201.500 90.200 ;
        RECT 203.800 87.900 204.200 90.200 ;
        RECT 1.400 70.800 1.800 73.100 ;
        RECT 4.100 70.800 4.600 72.100 ;
        RECT 5.800 70.800 6.200 72.100 ;
        RECT 8.600 70.800 9.000 73.000 ;
        RECT 10.200 70.800 10.600 72.100 ;
        RECT 11.800 70.800 12.200 72.100 ;
        RECT 12.600 70.800 13.000 72.100 ;
        RECT 14.700 70.800 15.100 73.100 ;
        RECT 17.400 70.800 17.800 72.700 ;
        RECT 19.800 70.800 20.200 73.100 ;
        RECT 22.500 70.800 23.000 72.100 ;
        RECT 24.200 70.800 24.600 72.100 ;
        RECT 27.000 70.800 27.400 73.000 ;
        RECT 28.600 70.800 29.000 73.100 ;
        RECT 31.800 70.800 32.200 72.100 ;
        RECT 33.400 70.800 33.800 73.100 ;
        RECT 36.100 70.800 36.600 72.100 ;
        RECT 37.800 70.800 38.200 72.100 ;
        RECT 40.600 70.800 41.000 73.000 ;
        RECT 42.200 70.800 42.600 73.100 ;
        RECT 46.200 70.800 46.600 72.700 ;
        RECT 48.600 70.800 49.000 72.700 ;
        RECT 53.400 70.800 53.800 72.700 ;
        RECT 55.800 70.800 56.200 73.100 ;
        RECT 57.400 70.800 57.800 73.100 ;
        RECT 59.000 70.800 59.400 72.100 ;
        RECT 60.600 70.800 61.000 72.100 ;
        RECT 63.800 70.800 64.200 72.700 ;
        RECT 66.200 70.800 66.600 72.700 ;
        RECT 69.400 70.800 69.800 72.700 ;
        RECT 74.200 70.800 74.600 72.700 ;
        RECT 78.200 70.800 78.600 72.700 ;
        RECT 82.200 70.800 82.600 72.700 ;
        RECT 84.600 70.800 85.000 72.700 ;
        RECT 87.000 70.800 87.400 72.100 ;
        RECT 89.100 70.800 89.500 73.100 ;
        RECT 91.000 70.800 91.400 72.700 ;
        RECT 94.200 70.800 94.600 72.100 ;
        RECT 95.800 70.800 96.200 72.100 ;
        RECT 97.400 70.800 97.800 73.000 ;
        RECT 100.200 70.800 100.600 72.100 ;
        RECT 101.800 70.800 102.300 72.100 ;
        RECT 104.600 70.800 105.000 73.100 ;
        RECT 107.800 70.800 108.200 73.100 ;
        RECT 111.800 70.800 112.200 72.700 ;
        RECT 113.400 70.800 113.800 72.100 ;
        RECT 115.000 70.800 115.400 72.100 ;
        RECT 117.400 70.800 117.800 72.700 ;
        RECT 119.800 70.800 120.200 73.000 ;
        RECT 122.600 70.800 123.000 72.100 ;
        RECT 124.200 70.800 124.700 72.100 ;
        RECT 127.000 70.800 127.400 73.100 ;
        RECT 128.600 70.800 129.000 72.100 ;
        RECT 130.200 70.800 130.600 72.100 ;
        RECT 131.000 70.800 131.400 72.100 ;
        RECT 132.600 70.800 133.000 72.100 ;
        RECT 133.400 70.800 133.800 72.100 ;
        RECT 135.500 70.800 135.900 73.100 ;
        RECT 137.400 70.800 137.800 72.700 ;
        RECT 141.400 70.800 141.800 73.100 ;
        RECT 143.000 70.800 143.400 73.100 ;
        RECT 145.700 70.800 146.200 72.100 ;
        RECT 147.400 70.800 147.800 72.100 ;
        RECT 150.200 70.800 150.600 73.000 ;
        RECT 153.700 70.800 154.100 73.100 ;
        RECT 155.800 70.800 156.200 72.100 ;
        RECT 156.600 70.800 157.000 72.100 ;
        RECT 159.800 70.800 160.200 72.700 ;
        RECT 163.000 70.800 163.400 73.100 ;
        RECT 163.800 70.800 164.200 72.100 ;
        RECT 165.400 70.800 165.800 72.100 ;
        RECT 166.200 70.800 166.600 72.100 ;
        RECT 168.300 70.800 168.700 73.100 ;
        RECT 170.200 70.800 170.600 73.100 ;
        RECT 171.800 70.800 172.200 73.100 ;
        RECT 172.600 70.800 173.000 72.100 ;
        RECT 174.700 70.800 175.100 73.100 ;
        RECT 175.800 70.800 176.200 72.100 ;
        RECT 177.400 70.800 177.800 72.100 ;
        RECT 178.200 70.800 178.600 72.100 ;
        RECT 180.300 70.800 180.700 73.100 ;
        RECT 182.200 70.800 182.600 73.000 ;
        RECT 185.000 70.800 185.400 72.100 ;
        RECT 186.600 70.800 187.100 72.100 ;
        RECT 189.400 70.800 189.800 73.100 ;
        RECT 191.800 70.800 192.200 72.100 ;
        RECT 192.900 70.800 193.300 73.100 ;
        RECT 195.000 70.800 195.400 72.100 ;
        RECT 196.600 70.800 197.000 73.000 ;
        RECT 199.400 70.800 199.800 72.100 ;
        RECT 201.000 70.800 201.500 72.100 ;
        RECT 203.800 70.800 204.200 73.100 ;
        RECT 0.200 70.200 205.400 70.800 ;
        RECT 1.400 67.900 1.800 70.200 ;
        RECT 4.100 68.900 4.600 70.200 ;
        RECT 5.800 68.900 6.200 70.200 ;
        RECT 8.600 68.000 9.000 70.200 ;
        RECT 11.800 68.300 12.200 70.200 ;
        RECT 15.000 67.900 15.400 70.200 ;
        RECT 16.600 67.900 17.000 70.200 ;
        RECT 19.300 68.900 19.800 70.200 ;
        RECT 21.000 68.900 21.400 70.200 ;
        RECT 23.800 68.000 24.200 70.200 ;
        RECT 26.200 68.300 26.600 70.200 ;
        RECT 29.400 68.300 29.800 70.200 ;
        RECT 33.400 67.900 33.800 70.200 ;
        RECT 35.000 67.900 35.400 70.200 ;
        RECT 37.700 68.900 38.200 70.200 ;
        RECT 39.400 68.900 39.800 70.200 ;
        RECT 42.200 68.000 42.600 70.200 ;
        RECT 44.600 68.300 45.000 70.200 ;
        RECT 47.300 67.900 47.700 70.200 ;
        RECT 49.400 68.900 49.800 70.200 ;
        RECT 52.600 68.300 53.000 70.200 ;
        RECT 56.600 68.300 57.000 70.200 ;
        RECT 59.800 67.900 60.200 70.200 ;
        RECT 61.400 67.900 61.800 70.200 ;
        RECT 64.100 68.900 64.600 70.200 ;
        RECT 65.800 68.900 66.200 70.200 ;
        RECT 68.600 68.000 69.000 70.200 ;
        RECT 70.500 67.900 70.900 70.200 ;
        RECT 72.600 68.900 73.000 70.200 ;
        RECT 73.400 68.900 73.800 70.200 ;
        RECT 75.000 68.900 75.400 70.200 ;
        RECT 76.600 67.900 77.000 70.200 ;
        RECT 78.200 67.900 78.600 70.200 ;
        RECT 80.600 67.900 81.000 70.200 ;
        RECT 83.000 68.300 83.400 70.200 ;
        RECT 86.200 68.300 86.600 70.200 ;
        RECT 89.400 67.900 89.800 70.200 ;
        RECT 91.800 68.300 92.200 70.200 ;
        RECT 95.000 67.900 95.400 70.200 ;
        RECT 97.400 68.300 97.800 70.200 ;
        RECT 99.000 68.900 99.400 70.200 ;
        RECT 101.100 67.900 101.500 70.200 ;
        RECT 105.400 68.300 105.800 70.200 ;
        RECT 107.800 67.900 108.200 70.200 ;
        RECT 110.500 68.900 111.000 70.200 ;
        RECT 112.200 68.900 112.600 70.200 ;
        RECT 115.000 68.000 115.400 70.200 ;
        RECT 116.900 67.900 117.300 70.200 ;
        RECT 119.000 68.900 119.400 70.200 ;
        RECT 120.600 68.000 121.000 70.200 ;
        RECT 123.400 68.900 123.800 70.200 ;
        RECT 125.000 68.900 125.500 70.200 ;
        RECT 127.800 67.900 128.200 70.200 ;
        RECT 129.400 68.900 129.800 70.200 ;
        RECT 131.500 67.900 131.900 70.200 ;
        RECT 132.600 67.900 133.000 70.200 ;
        RECT 136.600 68.300 137.000 70.200 ;
        RECT 138.500 67.900 138.900 70.200 ;
        RECT 140.600 68.900 141.000 70.200 ;
        RECT 142.200 67.900 142.600 70.200 ;
        RECT 143.800 67.900 144.200 70.200 ;
        RECT 146.200 68.300 146.600 70.200 ;
        RECT 148.100 67.900 148.500 70.200 ;
        RECT 150.200 68.900 150.600 70.200 ;
        RECT 151.800 68.300 152.200 70.200 ;
        RECT 156.600 67.900 157.000 70.200 ;
        RECT 159.300 68.900 159.800 70.200 ;
        RECT 161.000 68.900 161.400 70.200 ;
        RECT 163.800 68.000 164.200 70.200 ;
        RECT 166.200 67.700 166.600 70.200 ;
        RECT 168.800 67.500 169.200 70.200 ;
        RECT 171.000 68.900 171.400 70.200 ;
        RECT 172.600 68.000 173.000 70.200 ;
        RECT 175.400 68.900 175.800 70.200 ;
        RECT 177.000 68.900 177.500 70.200 ;
        RECT 179.800 67.900 180.200 70.200 ;
        RECT 182.000 67.500 182.400 70.200 ;
        RECT 184.600 67.700 185.000 70.200 ;
        RECT 186.500 67.900 186.900 70.200 ;
        RECT 188.600 68.900 189.000 70.200 ;
        RECT 191.000 68.300 191.400 70.200 ;
        RECT 192.600 67.900 193.000 70.200 ;
        RECT 194.200 67.900 194.600 70.200 ;
        RECT 196.600 68.300 197.000 70.200 ;
        RECT 198.200 68.900 198.600 70.200 ;
        RECT 199.800 68.900 200.200 70.200 ;
        RECT 200.600 68.900 201.000 70.200 ;
        RECT 202.700 67.900 203.100 70.200 ;
        RECT 1.400 50.800 1.800 53.100 ;
        RECT 4.100 50.800 4.600 52.100 ;
        RECT 5.800 50.800 6.200 52.100 ;
        RECT 8.600 50.800 9.000 53.000 ;
        RECT 11.000 50.800 11.400 53.100 ;
        RECT 13.700 50.800 14.200 52.100 ;
        RECT 15.400 50.800 15.800 52.100 ;
        RECT 18.200 50.800 18.600 53.000 ;
        RECT 20.600 50.800 21.000 52.700 ;
        RECT 24.600 50.800 25.000 53.100 ;
        RECT 26.200 50.800 26.600 53.100 ;
        RECT 28.900 50.800 29.400 52.100 ;
        RECT 30.600 50.800 31.000 52.100 ;
        RECT 33.400 50.800 33.800 53.000 ;
        RECT 35.000 50.800 35.400 53.100 ;
        RECT 39.000 50.800 39.400 52.700 ;
        RECT 41.400 50.800 41.800 52.700 ;
        RECT 44.600 50.800 45.000 53.100 ;
        RECT 47.300 50.800 47.800 52.100 ;
        RECT 49.000 50.800 49.400 52.100 ;
        RECT 51.800 50.800 52.200 53.000 ;
        RECT 55.800 50.800 56.200 52.700 ;
        RECT 59.800 50.800 60.200 53.100 ;
        RECT 62.200 50.800 62.600 52.700 ;
        RECT 64.100 50.800 64.500 53.100 ;
        RECT 66.200 50.800 66.600 52.100 ;
        RECT 67.800 50.800 68.200 53.100 ;
        RECT 70.500 50.800 71.000 52.100 ;
        RECT 72.200 50.800 72.600 52.100 ;
        RECT 75.000 50.800 75.400 53.000 ;
        RECT 77.400 50.800 77.800 52.700 ;
        RECT 81.400 50.800 81.800 53.100 ;
        RECT 82.200 50.800 82.600 52.100 ;
        RECT 84.300 50.800 84.700 53.100 ;
        RECT 87.000 50.800 87.400 52.700 ;
        RECT 89.400 50.800 89.800 52.700 ;
        RECT 93.400 50.800 93.800 53.100 ;
        RECT 95.000 50.800 95.400 53.100 ;
        RECT 97.700 50.800 98.200 52.100 ;
        RECT 99.400 50.800 99.800 52.100 ;
        RECT 102.200 50.800 102.600 53.000 ;
        RECT 107.000 50.800 107.400 52.700 ;
        RECT 109.400 50.800 109.800 52.100 ;
        RECT 110.200 50.800 110.600 53.100 ;
        RECT 114.200 50.800 114.600 52.700 ;
        RECT 116.100 50.800 116.500 53.100 ;
        RECT 118.200 50.800 118.600 52.100 ;
        RECT 119.800 50.800 120.200 53.000 ;
        RECT 122.600 50.800 123.000 52.100 ;
        RECT 124.200 50.800 124.700 52.100 ;
        RECT 127.000 50.800 127.400 53.100 ;
        RECT 129.400 50.800 129.800 52.700 ;
        RECT 133.400 50.800 133.800 53.100 ;
        RECT 135.000 50.800 135.400 53.100 ;
        RECT 137.700 50.800 138.200 52.100 ;
        RECT 139.400 50.800 139.800 52.100 ;
        RECT 142.200 50.800 142.600 53.000 ;
        RECT 144.600 50.800 145.000 53.100 ;
        RECT 146.200 50.800 146.600 53.100 ;
        RECT 147.800 50.800 148.200 53.000 ;
        RECT 150.600 50.800 151.000 52.100 ;
        RECT 152.200 50.800 152.700 52.100 ;
        RECT 155.000 50.800 155.400 53.100 ;
        RECT 159.000 50.800 159.400 52.100 ;
        RECT 160.600 50.800 161.000 53.000 ;
        RECT 163.400 50.800 163.800 52.100 ;
        RECT 165.000 50.800 165.500 52.100 ;
        RECT 167.800 50.800 168.200 53.100 ;
        RECT 170.200 50.800 170.600 53.300 ;
        RECT 172.800 50.800 173.200 53.500 ;
        RECT 174.500 50.800 174.900 53.100 ;
        RECT 176.600 50.800 177.000 52.100 ;
        RECT 179.000 50.800 179.400 52.700 ;
        RECT 181.400 50.800 181.800 53.100 ;
        RECT 184.100 50.800 184.600 52.100 ;
        RECT 185.800 50.800 186.200 52.100 ;
        RECT 188.600 50.800 189.000 53.000 ;
        RECT 190.200 50.800 190.600 52.100 ;
        RECT 193.400 50.800 193.800 53.100 ;
        RECT 194.500 50.800 194.900 53.100 ;
        RECT 196.600 50.800 197.000 52.100 ;
        RECT 197.400 50.800 197.800 52.100 ;
        RECT 199.000 50.800 199.400 52.100 ;
        RECT 201.400 50.800 201.800 53.100 ;
        RECT 202.200 50.800 202.600 52.100 ;
        RECT 204.300 50.800 204.700 53.100 ;
        RECT 0.200 50.200 205.400 50.800 ;
        RECT 0.600 47.900 1.000 50.200 ;
        RECT 2.200 47.900 2.600 50.200 ;
        RECT 3.800 47.900 4.200 50.200 ;
        RECT 5.400 47.900 5.800 50.200 ;
        RECT 7.000 47.900 7.400 50.200 ;
        RECT 7.800 48.900 8.200 50.200 ;
        RECT 9.400 48.900 9.800 50.200 ;
        RECT 10.200 48.900 10.600 50.200 ;
        RECT 12.300 47.900 12.700 50.200 ;
        RECT 13.400 47.900 13.800 50.200 ;
        RECT 17.400 48.300 17.800 50.200 ;
        RECT 19.800 48.300 20.200 50.200 ;
        RECT 23.800 47.900 24.200 50.200 ;
        RECT 25.400 47.900 25.800 50.200 ;
        RECT 28.100 48.900 28.600 50.200 ;
        RECT 29.800 48.900 30.200 50.200 ;
        RECT 32.600 48.000 33.000 50.200 ;
        RECT 35.000 48.300 35.400 50.200 ;
        RECT 39.000 47.900 39.400 50.200 ;
        RECT 40.600 47.900 41.000 50.200 ;
        RECT 43.300 48.900 43.800 50.200 ;
        RECT 45.000 48.900 45.400 50.200 ;
        RECT 47.800 48.000 48.200 50.200 ;
        RECT 51.800 48.300 52.200 50.200 ;
        RECT 55.000 48.300 55.400 50.200 ;
        RECT 58.200 47.900 58.600 50.200 ;
        RECT 59.800 47.900 60.200 50.200 ;
        RECT 61.400 47.900 61.800 50.200 ;
        RECT 64.100 48.900 64.600 50.200 ;
        RECT 65.800 48.900 66.200 50.200 ;
        RECT 68.600 48.000 69.000 50.200 ;
        RECT 71.000 47.900 71.400 50.200 ;
        RECT 73.700 48.900 74.200 50.200 ;
        RECT 75.400 48.900 75.800 50.200 ;
        RECT 78.200 48.000 78.600 50.200 ;
        RECT 79.800 48.900 80.200 50.200 ;
        RECT 82.000 47.500 82.400 50.200 ;
        RECT 84.600 47.700 85.000 50.200 ;
        RECT 86.200 48.900 86.600 50.200 ;
        RECT 87.800 48.900 88.200 50.200 ;
        RECT 88.900 47.900 89.300 50.200 ;
        RECT 91.000 48.900 91.400 50.200 ;
        RECT 92.600 48.300 93.000 50.200 ;
        RECT 96.600 48.300 97.000 50.200 ;
        RECT 99.000 47.900 99.400 50.200 ;
        RECT 100.600 47.900 101.000 50.200 ;
        RECT 103.300 47.900 103.700 50.200 ;
        RECT 105.400 48.900 105.800 50.200 ;
        RECT 106.500 47.900 106.900 50.200 ;
        RECT 108.600 48.900 109.000 50.200 ;
        RECT 109.400 48.900 109.800 50.200 ;
        RECT 111.500 47.900 111.900 50.200 ;
        RECT 114.200 48.300 114.600 50.200 ;
        RECT 115.800 48.900 116.200 50.200 ;
        RECT 117.400 48.900 117.800 50.200 ;
        RECT 119.000 48.000 119.400 50.200 ;
        RECT 121.800 48.900 122.200 50.200 ;
        RECT 123.400 48.900 123.900 50.200 ;
        RECT 126.200 47.900 126.600 50.200 ;
        RECT 129.400 48.300 129.800 50.200 ;
        RECT 131.000 47.900 131.400 50.200 ;
        RECT 132.600 47.900 133.000 50.200 ;
        RECT 135.000 48.000 135.400 50.200 ;
        RECT 137.800 48.900 138.200 50.200 ;
        RECT 139.400 48.900 139.900 50.200 ;
        RECT 142.200 47.900 142.600 50.200 ;
        RECT 143.800 48.900 144.200 50.200 ;
        RECT 145.400 48.900 145.800 50.200 ;
        RECT 146.200 48.900 146.600 50.200 ;
        RECT 148.300 47.900 148.700 50.200 ;
        RECT 151.000 48.300 151.400 50.200 ;
        RECT 154.200 47.900 154.600 50.200 ;
        RECT 155.800 47.900 156.200 50.200 ;
        RECT 157.400 47.700 157.800 50.200 ;
        RECT 160.000 47.500 160.400 50.200 ;
        RECT 161.700 47.900 162.100 50.200 ;
        RECT 163.800 48.900 164.200 50.200 ;
        RECT 166.200 48.300 166.600 50.200 ;
        RECT 167.800 47.900 168.200 50.200 ;
        RECT 171.800 47.900 172.200 50.200 ;
        RECT 172.600 47.900 173.000 50.200 ;
        RECT 174.200 47.900 174.600 50.200 ;
        RECT 175.800 47.900 176.200 50.200 ;
        RECT 178.500 48.900 179.000 50.200 ;
        RECT 180.200 48.900 180.600 50.200 ;
        RECT 183.000 48.000 183.400 50.200 ;
        RECT 184.600 48.900 185.000 50.200 ;
        RECT 187.000 47.700 187.400 50.200 ;
        RECT 189.600 47.500 190.000 50.200 ;
        RECT 191.800 47.900 192.200 50.200 ;
        RECT 194.500 48.900 195.000 50.200 ;
        RECT 196.200 48.900 196.600 50.200 ;
        RECT 199.000 48.000 199.400 50.200 ;
        RECT 200.600 47.900 201.000 50.200 ;
        RECT 202.200 47.900 202.600 50.200 ;
        RECT 203.000 48.900 203.400 50.200 ;
        RECT 204.600 48.900 205.000 50.200 ;
        RECT 0.600 30.800 1.000 32.100 ;
        RECT 3.000 30.800 3.400 33.100 ;
        RECT 5.700 30.800 6.200 32.100 ;
        RECT 7.400 30.800 7.800 32.100 ;
        RECT 10.200 30.800 10.600 33.000 ;
        RECT 12.400 30.800 12.800 33.500 ;
        RECT 15.000 30.800 15.400 33.300 ;
        RECT 16.600 30.800 17.000 32.100 ;
        RECT 19.000 30.800 19.400 33.300 ;
        RECT 21.600 30.800 22.000 33.500 ;
        RECT 23.800 30.800 24.200 33.100 ;
        RECT 26.500 30.800 27.000 32.100 ;
        RECT 28.200 30.800 28.600 32.100 ;
        RECT 31.000 30.800 31.400 33.000 ;
        RECT 33.400 30.800 33.800 32.700 ;
        RECT 35.800 30.800 36.200 33.100 ;
        RECT 38.200 30.800 38.600 32.100 ;
        RECT 40.100 30.800 40.500 33.100 ;
        RECT 42.200 30.800 42.600 32.100 ;
        RECT 43.800 30.800 44.200 32.700 ;
        RECT 46.500 30.800 46.900 33.100 ;
        RECT 48.600 30.800 49.000 32.100 ;
        RECT 51.300 30.800 51.700 33.100 ;
        RECT 53.400 30.800 53.800 32.100 ;
        RECT 54.200 30.800 54.600 32.100 ;
        RECT 55.800 30.800 56.200 32.100 ;
        RECT 56.600 30.800 57.000 32.100 ;
        RECT 58.200 30.800 58.600 32.100 ;
        RECT 60.600 30.800 61.000 32.700 ;
        RECT 62.200 30.800 62.600 33.100 ;
        RECT 63.800 30.800 64.200 33.100 ;
        RECT 66.200 30.800 66.600 32.700 ;
        RECT 70.200 30.800 70.600 33.100 ;
        RECT 71.000 30.800 71.400 33.100 ;
        RECT 72.600 30.800 73.000 33.100 ;
        RECT 74.200 30.800 74.600 33.100 ;
        RECT 75.800 30.800 76.200 33.100 ;
        RECT 77.400 30.800 77.800 33.100 ;
        RECT 78.200 30.800 78.600 32.100 ;
        RECT 79.800 30.800 80.200 32.100 ;
        RECT 82.200 30.800 82.600 32.700 ;
        RECT 84.600 30.800 85.000 32.700 ;
        RECT 88.600 30.800 89.000 33.100 ;
        RECT 90.200 30.800 90.600 33.000 ;
        RECT 93.000 30.800 93.400 32.100 ;
        RECT 94.600 30.800 95.100 32.100 ;
        RECT 97.400 30.800 97.800 33.100 ;
        RECT 99.000 30.800 99.400 32.100 ;
        RECT 100.600 30.800 101.000 32.100 ;
        RECT 103.800 30.800 104.200 32.700 ;
        RECT 107.600 30.800 108.000 33.500 ;
        RECT 110.200 30.800 110.600 33.300 ;
        RECT 112.100 30.800 112.500 33.100 ;
        RECT 114.200 30.800 114.600 32.100 ;
        RECT 115.800 30.800 116.200 32.100 ;
        RECT 117.400 30.800 117.800 33.000 ;
        RECT 120.200 30.800 120.600 32.100 ;
        RECT 121.800 30.800 122.300 32.100 ;
        RECT 124.600 30.800 125.000 33.100 ;
        RECT 126.200 30.800 126.600 32.100 ;
        RECT 127.800 30.800 128.200 32.100 ;
        RECT 128.600 30.800 129.000 32.100 ;
        RECT 130.700 30.800 131.100 33.100 ;
        RECT 132.400 30.800 132.800 33.500 ;
        RECT 135.000 30.800 135.400 33.300 ;
        RECT 137.400 30.800 137.800 32.100 ;
        RECT 139.000 30.800 139.400 33.000 ;
        RECT 141.800 30.800 142.200 32.100 ;
        RECT 143.400 30.800 143.900 32.100 ;
        RECT 146.200 30.800 146.600 33.100 ;
        RECT 147.800 30.800 148.200 33.100 ;
        RECT 149.400 30.800 149.800 33.100 ;
        RECT 151.000 30.800 151.400 33.100 ;
        RECT 152.600 30.800 153.000 33.100 ;
        RECT 154.200 30.800 154.600 33.100 ;
        RECT 157.400 30.800 157.800 32.100 ;
        RECT 159.000 30.800 159.400 33.000 ;
        RECT 161.800 30.800 162.200 32.100 ;
        RECT 163.400 30.800 163.900 32.100 ;
        RECT 166.200 30.800 166.600 33.100 ;
        RECT 167.800 30.800 168.200 32.100 ;
        RECT 169.400 30.800 169.800 32.100 ;
        RECT 170.200 30.800 170.600 32.100 ;
        RECT 172.300 30.800 172.700 33.100 ;
        RECT 174.200 30.800 174.600 33.300 ;
        RECT 176.800 30.800 177.200 33.500 ;
        RECT 179.000 30.800 179.400 32.100 ;
        RECT 179.800 30.800 180.200 32.100 ;
        RECT 181.400 30.800 181.800 32.100 ;
        RECT 182.200 30.800 182.600 32.100 ;
        RECT 184.300 30.800 184.700 33.100 ;
        RECT 186.200 30.800 186.600 33.000 ;
        RECT 189.000 30.800 189.400 32.100 ;
        RECT 190.600 30.800 191.100 32.100 ;
        RECT 193.400 30.800 193.800 33.100 ;
        RECT 195.800 30.800 196.200 33.000 ;
        RECT 198.600 30.800 199.000 32.100 ;
        RECT 200.200 30.800 200.700 32.100 ;
        RECT 203.000 30.800 203.400 33.100 ;
        RECT 0.200 30.200 205.400 30.800 ;
        RECT 1.400 28.000 1.800 30.200 ;
        RECT 4.200 28.900 4.600 30.200 ;
        RECT 5.800 28.900 6.300 30.200 ;
        RECT 8.600 27.900 9.000 30.200 ;
        RECT 11.000 28.000 11.400 30.200 ;
        RECT 13.800 28.900 14.200 30.200 ;
        RECT 15.400 28.900 15.900 30.200 ;
        RECT 18.200 27.900 18.600 30.200 ;
        RECT 20.600 27.900 21.000 30.200 ;
        RECT 23.300 28.900 23.800 30.200 ;
        RECT 25.000 28.900 25.400 30.200 ;
        RECT 27.800 28.000 28.200 30.200 ;
        RECT 29.400 27.900 29.800 30.200 ;
        RECT 33.400 28.300 33.800 30.200 ;
        RECT 35.800 27.900 36.200 30.200 ;
        RECT 38.500 28.900 39.000 30.200 ;
        RECT 40.200 28.900 40.600 30.200 ;
        RECT 43.000 28.000 43.400 30.200 ;
        RECT 45.400 28.300 45.800 30.200 ;
        RECT 49.400 27.900 49.800 30.200 ;
        RECT 51.800 27.900 52.200 30.200 ;
        RECT 53.400 27.900 53.800 30.200 ;
        RECT 55.800 28.300 56.200 30.200 ;
        RECT 58.200 28.900 58.600 30.200 ;
        RECT 60.300 27.900 60.700 30.200 ;
        RECT 61.400 28.900 61.800 30.200 ;
        RECT 63.000 28.900 63.400 30.200 ;
        RECT 65.400 28.300 65.800 30.200 ;
        RECT 67.800 28.300 68.200 30.200 ;
        RECT 71.800 28.300 72.200 30.200 ;
        RECT 74.000 27.500 74.400 30.200 ;
        RECT 76.600 27.700 77.000 30.200 ;
        RECT 78.200 27.900 78.600 30.200 ;
        RECT 82.200 28.300 82.600 30.200 ;
        RECT 84.600 28.300 85.000 30.200 ;
        RECT 87.800 27.700 88.200 30.200 ;
        RECT 90.400 27.500 90.800 30.200 ;
        RECT 92.600 28.300 93.000 30.200 ;
        RECT 95.800 28.300 96.200 30.200 ;
        RECT 99.000 27.700 99.400 30.200 ;
        RECT 101.600 27.500 102.000 30.200 ;
        RECT 104.600 28.900 105.000 30.200 ;
        RECT 106.700 27.900 107.100 30.200 ;
        RECT 107.800 28.900 108.200 30.200 ;
        RECT 109.400 28.900 109.800 30.200 ;
        RECT 110.200 28.900 110.600 30.200 ;
        RECT 112.300 27.900 112.700 30.200 ;
        RECT 115.000 28.300 115.400 30.200 ;
        RECT 118.200 28.300 118.600 30.200 ;
        RECT 121.400 28.300 121.800 30.200 ;
        RECT 123.800 28.300 124.200 30.200 ;
        RECT 126.500 27.900 126.900 30.200 ;
        RECT 128.600 28.900 129.000 30.200 ;
        RECT 131.000 28.300 131.400 30.200 ;
        RECT 133.400 28.000 133.800 30.200 ;
        RECT 136.200 28.900 136.600 30.200 ;
        RECT 137.800 28.900 138.300 30.200 ;
        RECT 140.600 27.900 141.000 30.200 ;
        RECT 142.200 28.900 142.600 30.200 ;
        RECT 143.800 28.900 144.200 30.200 ;
        RECT 145.400 28.000 145.800 30.200 ;
        RECT 148.200 28.900 148.600 30.200 ;
        RECT 149.800 28.900 150.300 30.200 ;
        RECT 152.600 27.900 153.000 30.200 ;
        RECT 156.100 27.900 156.500 30.200 ;
        RECT 158.200 28.900 158.600 30.200 ;
        RECT 159.000 28.900 159.400 30.200 ;
        RECT 160.600 28.900 161.000 30.200 ;
        RECT 161.400 28.900 161.800 30.200 ;
        RECT 163.500 27.900 163.900 30.200 ;
        RECT 166.200 28.300 166.600 30.200 ;
        RECT 168.600 28.000 169.000 30.200 ;
        RECT 171.400 28.900 171.800 30.200 ;
        RECT 173.000 28.900 173.500 30.200 ;
        RECT 175.800 27.900 176.200 30.200 ;
        RECT 178.200 28.000 178.600 30.200 ;
        RECT 181.000 28.900 181.400 30.200 ;
        RECT 182.600 28.900 183.100 30.200 ;
        RECT 185.400 27.900 185.800 30.200 ;
        RECT 187.800 27.700 188.200 30.200 ;
        RECT 190.400 27.500 190.800 30.200 ;
        RECT 192.600 27.900 193.000 30.200 ;
        RECT 194.200 28.900 194.600 30.200 ;
        RECT 195.800 27.700 196.200 30.200 ;
        RECT 198.400 27.500 198.800 30.200 ;
        RECT 200.600 27.900 201.000 30.200 ;
        RECT 203.000 27.900 203.400 30.200 ;
        RECT 1.400 10.800 1.800 13.100 ;
        RECT 4.100 10.800 4.600 12.100 ;
        RECT 5.800 10.800 6.200 12.100 ;
        RECT 8.600 10.800 9.000 13.000 ;
        RECT 10.500 10.800 10.900 13.100 ;
        RECT 12.600 10.800 13.000 12.100 ;
        RECT 13.400 10.800 13.800 12.100 ;
        RECT 15.000 10.800 15.400 12.100 ;
        RECT 16.600 10.800 17.000 13.100 ;
        RECT 19.300 10.800 19.800 12.100 ;
        RECT 21.000 10.800 21.400 12.100 ;
        RECT 23.800 10.800 24.200 13.000 ;
        RECT 26.200 10.800 26.600 12.700 ;
        RECT 30.200 10.800 30.600 13.100 ;
        RECT 31.800 10.800 32.200 12.700 ;
        RECT 35.800 10.800 36.200 13.100 ;
        RECT 36.600 10.800 37.000 12.100 ;
        RECT 38.200 10.800 38.600 13.100 ;
        RECT 41.400 10.800 41.800 13.100 ;
        RECT 44.100 10.800 44.600 12.100 ;
        RECT 45.800 10.800 46.200 12.100 ;
        RECT 48.600 10.800 49.000 13.000 ;
        RECT 52.600 10.800 53.000 12.700 ;
        RECT 56.600 10.800 57.000 13.100 ;
        RECT 57.400 10.800 57.800 12.100 ;
        RECT 59.000 10.800 59.400 12.100 ;
        RECT 59.800 10.800 60.200 12.100 ;
        RECT 61.400 10.800 61.800 12.100 ;
        RECT 63.000 10.800 63.400 13.000 ;
        RECT 65.800 10.800 66.200 12.100 ;
        RECT 67.400 10.800 67.900 12.100 ;
        RECT 70.200 10.800 70.600 13.100 ;
        RECT 72.600 10.800 73.000 12.700 ;
        RECT 75.800 10.800 76.200 12.700 ;
        RECT 80.600 10.800 81.000 12.700 ;
        RECT 82.200 10.800 82.600 12.100 ;
        RECT 83.800 10.800 84.200 13.100 ;
        RECT 87.800 10.800 88.200 12.700 ;
        RECT 90.200 10.800 90.600 13.100 ;
        RECT 92.900 10.800 93.400 12.100 ;
        RECT 94.600 10.800 95.000 12.100 ;
        RECT 97.400 10.800 97.800 13.000 ;
        RECT 99.800 10.800 100.200 12.100 ;
        RECT 100.600 10.800 101.000 12.100 ;
        RECT 102.200 10.800 102.600 12.100 ;
        RECT 105.400 10.800 105.800 13.000 ;
        RECT 108.200 10.800 108.600 12.100 ;
        RECT 109.800 10.800 110.300 12.100 ;
        RECT 112.600 10.800 113.000 13.100 ;
        RECT 114.200 10.800 114.600 13.100 ;
        RECT 118.200 10.800 118.600 12.700 ;
        RECT 120.600 10.800 121.000 13.100 ;
        RECT 123.300 10.800 123.800 12.100 ;
        RECT 125.000 10.800 125.400 12.100 ;
        RECT 127.800 10.800 128.200 13.000 ;
        RECT 129.400 10.800 129.800 13.100 ;
        RECT 131.000 10.800 131.400 13.100 ;
        RECT 132.600 10.800 133.000 13.100 ;
        RECT 134.200 10.800 134.600 13.100 ;
        RECT 135.800 10.800 136.200 13.100 ;
        RECT 137.400 10.800 137.800 13.300 ;
        RECT 140.000 10.800 140.400 13.500 ;
        RECT 141.400 10.800 141.800 12.100 ;
        RECT 143.000 10.800 143.400 12.100 ;
        RECT 143.800 10.800 144.200 12.100 ;
        RECT 145.900 10.800 146.300 13.100 ;
        RECT 147.800 10.800 148.200 13.000 ;
        RECT 150.600 10.800 151.000 12.100 ;
        RECT 152.200 10.800 152.700 12.100 ;
        RECT 155.000 10.800 155.400 13.100 ;
        RECT 158.200 10.800 158.600 12.100 ;
        RECT 159.800 10.800 160.200 12.100 ;
        RECT 160.600 10.800 161.000 12.100 ;
        RECT 162.700 10.800 163.100 13.100 ;
        RECT 163.800 10.800 164.200 12.100 ;
        RECT 165.400 10.800 165.800 12.100 ;
        RECT 166.200 10.800 166.600 12.100 ;
        RECT 168.300 10.800 168.700 13.100 ;
        RECT 169.400 10.800 169.800 13.100 ;
        RECT 171.000 10.800 171.400 13.100 ;
        RECT 172.600 10.800 173.000 13.100 ;
        RECT 174.200 10.800 174.600 13.100 ;
        RECT 175.800 10.800 176.200 13.100 ;
        RECT 176.600 10.800 177.000 12.100 ;
        RECT 178.200 10.800 178.600 12.100 ;
        RECT 179.000 10.800 179.400 12.100 ;
        RECT 181.100 10.800 181.500 13.100 ;
        RECT 182.200 10.800 182.600 12.100 ;
        RECT 183.800 10.800 184.200 12.100 ;
        RECT 184.600 10.800 185.000 12.100 ;
        RECT 186.700 10.800 187.100 13.100 ;
        RECT 188.600 10.800 189.000 13.100 ;
        RECT 191.300 10.800 191.800 12.100 ;
        RECT 193.000 10.800 193.400 12.100 ;
        RECT 195.800 10.800 196.200 13.000 ;
        RECT 198.200 10.800 198.600 13.100 ;
        RECT 200.600 10.800 201.000 12.100 ;
        RECT 202.200 10.800 202.600 13.100 ;
        RECT 0.200 10.200 205.400 10.800 ;
        RECT 0.600 7.900 1.000 10.200 ;
        RECT 2.200 7.900 2.600 10.200 ;
        RECT 3.800 7.900 4.200 10.200 ;
        RECT 5.400 7.900 5.800 10.200 ;
        RECT 7.000 7.900 7.400 10.200 ;
        RECT 7.800 7.900 8.200 10.200 ;
        RECT 9.400 7.900 9.800 10.200 ;
        RECT 11.000 7.900 11.400 10.200 ;
        RECT 12.600 7.900 13.000 10.200 ;
        RECT 14.200 7.900 14.600 10.200 ;
        RECT 15.800 7.900 16.200 10.200 ;
        RECT 18.500 8.900 19.000 10.200 ;
        RECT 20.200 8.900 20.600 10.200 ;
        RECT 23.000 8.000 23.400 10.200 ;
        RECT 24.600 8.900 25.000 10.200 ;
        RECT 26.200 8.900 26.600 10.200 ;
        RECT 27.000 8.900 27.400 10.200 ;
        RECT 29.100 7.900 29.500 10.200 ;
        RECT 31.000 7.900 31.400 10.200 ;
        RECT 33.700 8.900 34.200 10.200 ;
        RECT 35.400 8.900 35.800 10.200 ;
        RECT 38.200 8.000 38.600 10.200 ;
        RECT 41.400 8.300 41.800 10.200 ;
        RECT 43.800 8.000 44.200 10.200 ;
        RECT 46.600 8.900 47.000 10.200 ;
        RECT 48.200 8.900 48.700 10.200 ;
        RECT 51.000 7.900 51.400 10.200 ;
        RECT 55.000 7.900 55.400 10.200 ;
        RECT 57.700 8.900 58.200 10.200 ;
        RECT 59.400 8.900 59.800 10.200 ;
        RECT 62.200 8.000 62.600 10.200 ;
        RECT 63.800 7.900 64.200 10.200 ;
        RECT 67.800 8.300 68.200 10.200 ;
        RECT 70.200 7.900 70.600 10.200 ;
        RECT 72.900 8.900 73.400 10.200 ;
        RECT 74.600 8.900 75.000 10.200 ;
        RECT 77.400 8.000 77.800 10.200 ;
        RECT 80.600 7.900 81.000 10.200 ;
        RECT 82.200 8.000 82.600 10.200 ;
        RECT 85.000 8.900 85.400 10.200 ;
        RECT 86.600 8.900 87.100 10.200 ;
        RECT 89.400 7.900 89.800 10.200 ;
        RECT 91.800 8.000 92.200 10.200 ;
        RECT 94.600 8.900 95.000 10.200 ;
        RECT 96.200 8.900 96.700 10.200 ;
        RECT 99.000 7.900 99.400 10.200 ;
        RECT 103.000 8.000 103.400 10.200 ;
        RECT 105.800 8.900 106.200 10.200 ;
        RECT 107.400 8.900 107.900 10.200 ;
        RECT 110.200 7.900 110.600 10.200 ;
        RECT 111.800 7.900 112.200 10.200 ;
        RECT 115.800 8.300 116.200 10.200 ;
        RECT 117.400 8.900 117.800 10.200 ;
        RECT 119.000 8.900 119.400 10.200 ;
        RECT 119.800 8.900 120.200 10.200 ;
        RECT 121.900 7.900 122.300 10.200 ;
        RECT 123.800 8.000 124.200 10.200 ;
        RECT 126.600 8.900 127.000 10.200 ;
        RECT 128.200 8.900 128.700 10.200 ;
        RECT 131.000 7.900 131.400 10.200 ;
        RECT 133.400 8.900 133.800 10.200 ;
        RECT 135.000 8.000 135.400 10.200 ;
        RECT 137.800 8.900 138.200 10.200 ;
        RECT 139.400 8.900 139.900 10.200 ;
        RECT 142.200 7.900 142.600 10.200 ;
        RECT 143.800 7.900 144.200 10.200 ;
        RECT 145.400 7.900 145.800 10.200 ;
        RECT 147.000 7.900 147.400 10.200 ;
        RECT 148.600 7.900 149.000 10.200 ;
        RECT 150.200 7.900 150.600 10.200 ;
        RECT 153.400 8.000 153.800 10.200 ;
        RECT 156.200 8.900 156.600 10.200 ;
        RECT 157.800 8.900 158.300 10.200 ;
        RECT 160.600 7.900 161.000 10.200 ;
        RECT 162.200 8.900 162.600 10.200 ;
        RECT 164.600 8.000 165.000 10.200 ;
        RECT 167.400 8.900 167.800 10.200 ;
        RECT 169.000 8.900 169.500 10.200 ;
        RECT 171.800 7.900 172.200 10.200 ;
        RECT 174.200 8.000 174.600 10.200 ;
        RECT 177.000 8.900 177.400 10.200 ;
        RECT 178.600 8.900 179.100 10.200 ;
        RECT 181.400 7.900 181.800 10.200 ;
        RECT 183.800 8.000 184.200 10.200 ;
        RECT 186.600 8.900 187.000 10.200 ;
        RECT 188.200 8.900 188.700 10.200 ;
        RECT 191.000 7.900 191.400 10.200 ;
        RECT 193.400 7.900 193.800 10.200 ;
        RECT 196.100 8.900 196.600 10.200 ;
        RECT 197.800 8.900 198.200 10.200 ;
        RECT 200.600 8.000 201.000 10.200 ;
        RECT 202.200 7.900 202.600 10.200 ;
        RECT 203.800 7.900 204.200 10.200 ;
      LAYER via1 ;
        RECT 101.800 170.300 102.200 170.700 ;
        RECT 102.500 170.300 102.900 170.700 ;
        RECT 101.800 150.300 102.200 150.700 ;
        RECT 102.500 150.300 102.900 150.700 ;
        RECT 101.800 130.300 102.200 130.700 ;
        RECT 102.500 130.300 102.900 130.700 ;
        RECT 101.800 110.300 102.200 110.700 ;
        RECT 102.500 110.300 102.900 110.700 ;
        RECT 101.800 90.300 102.200 90.700 ;
        RECT 102.500 90.300 102.900 90.700 ;
        RECT 101.800 70.300 102.200 70.700 ;
        RECT 102.500 70.300 102.900 70.700 ;
        RECT 101.800 50.300 102.200 50.700 ;
        RECT 102.500 50.300 102.900 50.700 ;
        RECT 101.800 30.300 102.200 30.700 ;
        RECT 102.500 30.300 102.900 30.700 ;
        RECT 101.800 10.300 102.200 10.700 ;
        RECT 102.500 10.300 102.900 10.700 ;
      LAYER metal2 ;
        RECT 101.600 170.300 103.200 170.700 ;
        RECT 101.600 150.300 103.200 150.700 ;
        RECT 101.600 130.300 103.200 130.700 ;
        RECT 101.600 110.300 103.200 110.700 ;
        RECT 101.600 90.300 103.200 90.700 ;
        RECT 101.600 70.300 103.200 70.700 ;
        RECT 101.600 50.300 103.200 50.700 ;
        RECT 101.600 30.300 103.200 30.700 ;
        RECT 101.600 10.300 103.200 10.700 ;
      LAYER via2 ;
        RECT 101.800 170.300 102.200 170.700 ;
        RECT 102.500 170.300 102.900 170.700 ;
        RECT 101.800 150.300 102.200 150.700 ;
        RECT 102.500 150.300 102.900 150.700 ;
        RECT 101.800 130.300 102.200 130.700 ;
        RECT 102.500 130.300 102.900 130.700 ;
        RECT 101.800 110.300 102.200 110.700 ;
        RECT 102.500 110.300 102.900 110.700 ;
        RECT 101.800 90.300 102.200 90.700 ;
        RECT 102.500 90.300 102.900 90.700 ;
        RECT 101.800 70.300 102.200 70.700 ;
        RECT 102.500 70.300 102.900 70.700 ;
        RECT 101.800 50.300 102.200 50.700 ;
        RECT 102.500 50.300 102.900 50.700 ;
        RECT 101.800 30.300 102.200 30.700 ;
        RECT 102.500 30.300 102.900 30.700 ;
        RECT 101.800 10.300 102.200 10.700 ;
        RECT 102.500 10.300 102.900 10.700 ;
      LAYER metal3 ;
        RECT 101.600 170.300 103.200 170.700 ;
        RECT 101.600 150.300 103.200 150.700 ;
        RECT 101.600 130.300 103.200 130.700 ;
        RECT 101.600 110.300 103.200 110.700 ;
        RECT 101.600 90.300 103.200 90.700 ;
        RECT 101.600 70.300 103.200 70.700 ;
        RECT 101.600 50.300 103.200 50.700 ;
        RECT 101.600 30.300 103.200 30.700 ;
        RECT 101.600 10.300 103.200 10.700 ;
      LAYER via3 ;
        RECT 101.800 170.300 102.200 170.700 ;
        RECT 102.600 170.300 103.000 170.700 ;
        RECT 101.800 150.300 102.200 150.700 ;
        RECT 102.600 150.300 103.000 150.700 ;
        RECT 101.800 130.300 102.200 130.700 ;
        RECT 102.600 130.300 103.000 130.700 ;
        RECT 101.800 110.300 102.200 110.700 ;
        RECT 102.600 110.300 103.000 110.700 ;
        RECT 101.800 90.300 102.200 90.700 ;
        RECT 102.600 90.300 103.000 90.700 ;
        RECT 101.800 70.300 102.200 70.700 ;
        RECT 102.600 70.300 103.000 70.700 ;
        RECT 101.800 50.300 102.200 50.700 ;
        RECT 102.600 50.300 103.000 50.700 ;
        RECT 101.800 30.300 102.200 30.700 ;
        RECT 102.600 30.300 103.000 30.700 ;
        RECT 101.800 10.300 102.200 10.700 ;
        RECT 102.600 10.300 103.000 10.700 ;
      LAYER metal4 ;
        RECT 101.600 170.300 103.200 170.700 ;
        RECT 101.600 150.300 103.200 150.700 ;
        RECT 101.600 130.300 103.200 130.700 ;
        RECT 101.600 110.300 103.200 110.700 ;
        RECT 101.600 90.300 103.200 90.700 ;
        RECT 101.600 70.300 103.200 70.700 ;
        RECT 101.600 50.300 103.200 50.700 ;
        RECT 101.600 30.300 103.200 30.700 ;
        RECT 101.600 10.300 103.200 10.700 ;
      LAYER via4 ;
        RECT 101.800 170.300 102.200 170.700 ;
        RECT 102.500 170.300 102.900 170.700 ;
        RECT 101.800 150.300 102.200 150.700 ;
        RECT 102.500 150.300 102.900 150.700 ;
        RECT 101.800 130.300 102.200 130.700 ;
        RECT 102.500 130.300 102.900 130.700 ;
        RECT 101.800 110.300 102.200 110.700 ;
        RECT 102.500 110.300 102.900 110.700 ;
        RECT 101.800 90.300 102.200 90.700 ;
        RECT 102.500 90.300 102.900 90.700 ;
        RECT 101.800 70.300 102.200 70.700 ;
        RECT 102.500 70.300 102.900 70.700 ;
        RECT 101.800 50.300 102.200 50.700 ;
        RECT 102.500 50.300 102.900 50.700 ;
        RECT 101.800 30.300 102.200 30.700 ;
        RECT 102.500 30.300 102.900 30.700 ;
        RECT 101.800 10.300 102.200 10.700 ;
        RECT 102.500 10.300 102.900 10.700 ;
      LAYER metal5 ;
        RECT 101.600 170.200 103.200 170.700 ;
        RECT 101.600 150.200 103.200 150.700 ;
        RECT 101.600 130.200 103.200 130.700 ;
        RECT 101.600 110.200 103.200 110.700 ;
        RECT 101.600 90.200 103.200 90.700 ;
        RECT 101.600 70.200 103.200 70.700 ;
        RECT 101.600 50.200 103.200 50.700 ;
        RECT 101.600 30.200 103.200 30.700 ;
        RECT 101.600 10.200 103.200 10.700 ;
      LAYER via5 ;
        RECT 102.600 170.200 103.100 170.700 ;
        RECT 102.600 150.200 103.100 150.700 ;
        RECT 102.600 130.200 103.100 130.700 ;
        RECT 102.600 110.200 103.100 110.700 ;
        RECT 102.600 90.200 103.100 90.700 ;
        RECT 102.600 70.200 103.100 70.700 ;
        RECT 102.600 50.200 103.100 50.700 ;
        RECT 102.600 30.200 103.100 30.700 ;
        RECT 102.600 10.200 103.100 10.700 ;
      LAYER metal6 ;
        RECT 101.600 -3.000 103.200 183.000 ;
    END
  END gnd
  PIN clk
    PORT
      LAYER metal1 ;
        RECT 5.400 174.100 6.300 174.500 ;
        RECT 91.300 174.100 92.200 174.500 ;
        RECT 120.900 174.100 121.800 174.500 ;
        RECT 5.400 173.800 5.800 174.100 ;
        RECT 91.800 173.800 92.200 174.100 ;
        RECT 121.400 173.800 121.800 174.100 ;
        RECT 167.000 174.100 167.900 174.500 ;
        RECT 167.000 173.800 167.400 174.100 ;
        RECT 0.600 94.100 1.500 94.500 ;
        RECT 0.600 93.800 1.000 94.100 ;
        RECT 0.600 46.900 1.000 47.200 ;
        RECT 0.600 46.500 1.500 46.900 ;
        RECT 153.700 34.100 154.600 34.500 ;
        RECT 155.000 34.100 155.400 34.200 ;
        RECT 154.200 33.800 155.400 34.100 ;
        RECT 135.300 14.100 136.200 14.500 ;
        RECT 135.800 13.800 136.200 14.100 ;
        RECT 169.400 14.100 170.300 14.500 ;
        RECT 169.400 13.800 169.800 14.100 ;
        RECT 0.600 6.900 1.000 7.200 ;
        RECT 7.800 6.900 8.200 7.200 ;
        RECT 143.800 6.900 144.200 7.200 ;
        RECT 0.600 6.500 1.500 6.900 ;
        RECT 7.800 6.500 8.700 6.900 ;
        RECT 143.800 6.500 144.700 6.900 ;
      LAYER via1 ;
        RECT 0.600 46.800 1.000 47.200 ;
        RECT 155.000 33.800 155.400 34.200 ;
        RECT 0.600 6.800 1.000 7.200 ;
        RECT 7.800 6.800 8.200 7.200 ;
        RECT 143.800 6.800 144.200 7.200 ;
      LAYER metal2 ;
        RECT 11.800 182.800 12.200 183.200 ;
        RECT 11.800 179.200 12.100 182.800 ;
        RECT 5.400 178.800 5.800 179.200 ;
        RECT 11.800 178.800 12.200 179.200 ;
        RECT 91.800 178.800 92.200 179.200 ;
        RECT 5.400 174.200 5.700 178.800 ;
        RECT 91.800 175.200 92.100 178.800 ;
        RECT 91.800 174.800 92.200 175.200 ;
        RECT 121.400 174.800 121.800 175.200 ;
        RECT 91.800 174.200 92.100 174.800 ;
        RECT 121.400 174.200 121.700 174.800 ;
        RECT 5.400 173.800 5.800 174.200 ;
        RECT 91.800 173.800 92.200 174.200 ;
        RECT 121.400 173.800 121.800 174.200 ;
        RECT 166.200 174.100 166.600 174.200 ;
        RECT 167.000 174.100 167.400 174.200 ;
        RECT 166.200 173.800 167.400 174.100 ;
        RECT 5.400 159.200 5.700 173.800 ;
        RECT 5.400 158.800 5.800 159.200 ;
        RECT 0.600 98.800 1.000 99.200 ;
        RECT 0.600 94.200 0.900 98.800 ;
        RECT 0.600 93.800 1.000 94.200 ;
        RECT 0.600 47.100 1.000 47.200 ;
        RECT 1.400 47.100 1.800 47.200 ;
        RECT 0.600 46.800 1.800 47.100 ;
        RECT 155.000 33.800 155.400 34.200 ;
        RECT 155.000 15.200 155.300 33.800 ;
        RECT 135.800 14.800 136.200 15.200 ;
        RECT 143.800 14.800 144.200 15.200 ;
        RECT 155.000 14.800 155.400 15.200 ;
        RECT 169.400 14.800 169.800 15.200 ;
        RECT 135.800 14.200 136.100 14.800 ;
        RECT 135.800 13.800 136.200 14.200 ;
        RECT 143.800 7.200 144.100 14.800 ;
        RECT 169.400 14.200 169.700 14.800 ;
        RECT 169.400 13.800 169.800 14.200 ;
        RECT 0.600 7.100 1.000 7.200 ;
        RECT 1.400 7.100 1.800 7.200 ;
        RECT 0.600 6.800 1.800 7.100 ;
        RECT 7.000 7.100 7.400 7.200 ;
        RECT 7.800 7.100 8.200 7.200 ;
        RECT 7.000 6.800 8.200 7.100 ;
        RECT 143.800 6.800 144.200 7.200 ;
      LAYER via2 ;
        RECT 1.400 46.800 1.800 47.200 ;
        RECT 1.400 6.800 1.800 7.200 ;
      LAYER metal3 ;
        RECT 5.400 179.100 5.800 179.200 ;
        RECT 11.800 179.100 12.200 179.200 ;
        RECT 91.800 179.100 92.200 179.200 ;
        RECT 5.400 178.800 92.200 179.100 ;
        RECT 91.800 175.100 92.200 175.200 ;
        RECT 121.400 175.100 121.800 175.200 ;
        RECT 91.800 174.800 166.500 175.100 ;
        RECT 166.200 174.200 166.500 174.800 ;
        RECT 166.200 174.100 166.600 174.200 ;
        RECT 167.000 174.100 167.400 174.200 ;
        RECT 166.200 173.800 167.400 174.100 ;
        RECT 3.000 159.100 3.400 159.200 ;
        RECT 5.400 159.100 5.800 159.200 ;
        RECT 3.000 158.800 5.800 159.100 ;
        RECT 0.600 99.100 1.000 99.200 ;
        RECT 3.000 99.100 3.400 99.200 ;
        RECT 0.600 98.800 3.400 99.100 ;
        RECT 1.400 47.100 1.800 47.200 ;
        RECT 3.000 47.100 3.400 47.200 ;
        RECT 1.400 46.800 3.400 47.100 ;
        RECT 135.800 15.100 136.200 15.200 ;
        RECT 143.800 15.100 144.200 15.200 ;
        RECT 155.000 15.100 155.400 15.200 ;
        RECT 167.000 15.100 167.400 15.200 ;
        RECT 169.400 15.100 169.800 15.200 ;
        RECT 135.800 14.800 169.800 15.100 ;
        RECT 1.400 7.100 1.800 7.200 ;
        RECT 3.000 7.100 3.400 7.200 ;
        RECT 7.000 7.100 7.400 7.200 ;
        RECT 1.400 6.800 7.400 7.100 ;
      LAYER via3 ;
        RECT 167.000 173.800 167.400 174.200 ;
        RECT 3.000 98.800 3.400 99.200 ;
        RECT 3.000 46.800 3.400 47.200 ;
        RECT 167.000 14.800 167.400 15.200 ;
        RECT 3.000 6.800 3.400 7.200 ;
      LAYER metal4 ;
        RECT 167.000 173.800 167.400 174.200 ;
        RECT 3.000 158.800 3.400 159.200 ;
        RECT 3.000 99.200 3.300 158.800 ;
        RECT 3.000 98.800 3.400 99.200 ;
        RECT 3.000 47.200 3.300 98.800 ;
        RECT 3.000 46.800 3.400 47.200 ;
        RECT 3.000 7.200 3.300 46.800 ;
        RECT 167.000 15.200 167.300 173.800 ;
        RECT 167.000 14.800 167.400 15.200 ;
        RECT 3.000 6.800 3.400 7.200 ;
    END
  END clk
  PIN reset
    PORT
      LAYER metal1 ;
        RECT 81.400 173.400 81.800 174.200 ;
      LAYER via1 ;
        RECT 81.400 173.800 81.800 174.200 ;
      LAYER metal2 ;
        RECT 83.000 182.800 83.400 183.200 ;
        RECT 83.000 180.200 83.300 182.800 ;
        RECT 81.400 179.800 81.800 180.200 ;
        RECT 83.000 179.800 83.400 180.200 ;
        RECT 81.400 174.200 81.700 179.800 ;
        RECT 81.400 173.800 81.800 174.200 ;
      LAYER metal3 ;
        RECT 81.400 180.100 81.800 180.200 ;
        RECT 83.000 180.100 83.400 180.200 ;
        RECT 81.400 179.800 83.400 180.100 ;
    END
  END reset
  PIN d_in[0]
    PORT
      LAYER metal1 ;
        RECT 201.400 53.400 201.800 54.200 ;
        RECT 202.200 6.800 202.600 7.600 ;
      LAYER via1 ;
        RECT 201.400 53.800 201.800 54.200 ;
      LAYER metal2 ;
        RECT 201.400 53.800 201.800 54.200 ;
        RECT 201.400 51.200 201.700 53.800 ;
        RECT 201.400 50.800 201.800 51.200 ;
        RECT 202.200 6.800 202.600 7.200 ;
        RECT 202.200 6.200 202.500 6.800 ;
        RECT 202.200 5.800 202.600 6.200 ;
      LAYER metal3 ;
        RECT 201.400 51.100 201.800 51.200 ;
        RECT 204.600 51.100 205.000 51.200 ;
        RECT 201.400 50.800 205.000 51.100 ;
        RECT 202.200 6.100 202.600 6.200 ;
        RECT 204.600 6.100 205.000 6.200 ;
        RECT 207.800 6.100 208.200 6.200 ;
        RECT 202.200 5.800 208.200 6.100 ;
      LAYER via3 ;
        RECT 204.600 50.800 205.000 51.200 ;
        RECT 204.600 5.800 205.000 6.200 ;
      LAYER metal4 ;
        RECT 204.600 50.800 205.000 51.200 ;
        RECT 204.600 6.200 204.900 50.800 ;
        RECT 204.600 5.800 205.000 6.200 ;
    END
  END d_in[0]
  PIN d_in[1]
    PORT
      LAYER metal1 ;
        RECT 155.800 46.800 156.200 47.600 ;
        RECT 167.800 46.800 168.200 47.600 ;
      LAYER metal2 ;
        RECT 155.800 47.800 156.200 48.200 ;
        RECT 167.800 47.800 168.200 48.200 ;
        RECT 155.800 47.200 156.100 47.800 ;
        RECT 167.800 47.200 168.100 47.800 ;
        RECT 155.800 46.800 156.200 47.200 ;
        RECT 167.800 46.800 168.200 47.200 ;
        RECT 167.800 45.200 168.100 46.800 ;
        RECT 167.800 44.800 168.200 45.200 ;
      LAYER metal3 ;
        RECT 155.800 48.100 156.200 48.200 ;
        RECT 167.800 48.100 168.200 48.200 ;
        RECT 155.800 47.800 168.200 48.100 ;
        RECT 167.800 45.100 168.200 45.200 ;
        RECT 207.800 45.100 208.200 45.200 ;
        RECT 167.800 44.800 208.200 45.100 ;
    END
  END d_in[1]
  PIN d_in[2]
    PORT
      LAYER metal1 ;
        RECT 171.800 47.100 172.200 47.600 ;
        RECT 172.600 47.100 173.000 47.600 ;
        RECT 171.800 46.800 173.000 47.100 ;
      LAYER via1 ;
        RECT 172.600 46.800 173.000 47.200 ;
      LAYER metal2 ;
        RECT 172.600 48.800 173.000 49.200 ;
        RECT 172.600 47.200 172.900 48.800 ;
        RECT 172.600 46.800 173.000 47.200 ;
      LAYER metal3 ;
        RECT 172.600 49.100 173.000 49.200 ;
        RECT 203.800 49.100 204.200 49.200 ;
        RECT 172.600 48.800 204.200 49.100 ;
        RECT 203.800 47.100 204.200 47.200 ;
        RECT 207.800 47.100 208.200 47.200 ;
        RECT 203.800 46.800 208.200 47.100 ;
      LAYER via3 ;
        RECT 203.800 48.800 204.200 49.200 ;
      LAYER metal4 ;
        RECT 203.800 48.800 204.200 49.200 ;
        RECT 203.800 47.200 204.100 48.800 ;
        RECT 203.800 46.800 204.200 47.200 ;
    END
  END d_in[2]
  PIN d_in[3]
    PORT
      LAYER metal1 ;
        RECT 192.600 66.800 193.000 67.600 ;
        RECT 193.400 53.400 193.800 54.200 ;
      LAYER via1 ;
        RECT 193.400 53.800 193.800 54.200 ;
      LAYER metal2 ;
        RECT 192.600 66.800 193.000 67.200 ;
        RECT 192.600 66.200 192.900 66.800 ;
        RECT 192.600 65.800 193.000 66.200 ;
        RECT 192.600 54.100 193.000 54.200 ;
        RECT 193.400 54.100 193.800 54.200 ;
        RECT 192.600 53.800 193.800 54.100 ;
      LAYER metal3 ;
        RECT 192.600 66.100 193.000 66.200 ;
        RECT 193.400 66.100 193.800 66.200 ;
        RECT 192.600 65.800 193.800 66.100 ;
        RECT 207.800 54.800 208.200 55.200 ;
        RECT 192.600 54.100 193.000 54.200 ;
        RECT 193.400 54.100 193.800 54.200 ;
        RECT 207.800 54.100 208.100 54.800 ;
        RECT 192.600 53.800 208.100 54.100 ;
      LAYER via3 ;
        RECT 193.400 65.800 193.800 66.200 ;
        RECT 193.400 53.800 193.800 54.200 ;
      LAYER metal4 ;
        RECT 193.400 65.800 193.800 66.200 ;
        RECT 193.400 54.200 193.700 65.800 ;
        RECT 193.400 53.800 193.800 54.200 ;
    END
  END d_in[3]
  PIN d_in[4]
    PORT
      LAYER metal1 ;
        RECT 203.800 107.100 204.200 107.600 ;
        RECT 204.600 107.100 205.000 107.200 ;
        RECT 203.800 106.800 205.000 107.100 ;
        RECT 200.600 46.800 201.000 47.600 ;
      LAYER via1 ;
        RECT 204.600 106.800 205.000 107.200 ;
      LAYER metal2 ;
        RECT 204.600 106.800 205.000 107.200 ;
        RECT 204.600 105.200 204.900 106.800 ;
        RECT 204.600 104.800 205.000 105.200 ;
        RECT 200.600 51.800 201.000 52.200 ;
        RECT 200.600 47.200 200.900 51.800 ;
        RECT 200.600 46.800 201.000 47.200 ;
      LAYER metal3 ;
        RECT 203.800 105.100 204.200 105.200 ;
        RECT 204.600 105.100 205.000 105.200 ;
        RECT 207.800 105.100 208.200 105.200 ;
        RECT 203.800 104.800 208.200 105.100 ;
        RECT 200.600 52.100 201.000 52.200 ;
        RECT 203.800 52.100 204.200 52.200 ;
        RECT 200.600 51.800 204.200 52.100 ;
      LAYER via3 ;
        RECT 203.800 51.800 204.200 52.200 ;
      LAYER metal4 ;
        RECT 203.800 104.800 204.200 105.200 ;
        RECT 203.800 52.200 204.100 104.800 ;
        RECT 203.800 51.800 204.200 52.200 ;
    END
  END d_in[4]
  PIN d_in[5]
    PORT
      LAYER metal1 ;
        RECT 179.000 126.800 179.400 127.600 ;
        RECT 185.400 126.800 185.800 127.600 ;
      LAYER metal2 ;
        RECT 179.000 126.800 179.400 127.200 ;
        RECT 185.400 126.800 185.800 127.200 ;
        RECT 179.000 124.200 179.300 126.800 ;
        RECT 185.400 125.200 185.700 126.800 ;
        RECT 185.400 124.800 185.800 125.200 ;
        RECT 185.400 124.200 185.700 124.800 ;
        RECT 179.000 123.800 179.400 124.200 ;
        RECT 185.400 123.800 185.800 124.200 ;
      LAYER metal3 ;
        RECT 185.400 125.100 185.800 125.200 ;
        RECT 207.800 125.100 208.200 125.200 ;
        RECT 185.400 124.800 208.200 125.100 ;
        RECT 179.000 124.100 179.400 124.200 ;
        RECT 185.400 124.100 185.800 124.200 ;
        RECT 179.000 123.800 185.800 124.100 ;
    END
  END d_in[5]
  PIN d_in[6]
    PORT
      LAYER metal1 ;
        RECT 181.400 126.800 181.800 127.600 ;
        RECT 190.200 126.800 190.600 127.600 ;
      LAYER metal2 ;
        RECT 181.400 128.800 181.800 129.200 ;
        RECT 190.200 128.800 190.600 129.200 ;
        RECT 181.400 127.200 181.700 128.800 ;
        RECT 190.200 127.200 190.500 128.800 ;
        RECT 181.400 126.800 181.800 127.200 ;
        RECT 190.200 126.800 190.600 127.200 ;
      LAYER metal3 ;
        RECT 181.400 129.100 181.800 129.200 ;
        RECT 182.200 129.100 182.600 129.200 ;
        RECT 181.400 128.800 182.600 129.100 ;
        RECT 189.400 129.100 189.800 129.200 ;
        RECT 190.200 129.100 190.600 129.200 ;
        RECT 204.600 129.100 205.000 129.200 ;
        RECT 189.400 128.800 205.000 129.100 ;
        RECT 204.600 127.100 205.000 127.200 ;
        RECT 207.800 127.100 208.200 127.200 ;
        RECT 204.600 126.800 208.200 127.100 ;
      LAYER via3 ;
        RECT 182.200 128.800 182.600 129.200 ;
        RECT 204.600 128.800 205.000 129.200 ;
      LAYER metal4 ;
        RECT 182.200 129.100 182.600 129.200 ;
        RECT 183.000 129.100 183.400 129.200 ;
        RECT 182.200 128.800 183.400 129.100 ;
        RECT 188.600 129.100 189.000 129.200 ;
        RECT 189.400 129.100 189.800 129.200 ;
        RECT 188.600 128.800 189.800 129.100 ;
        RECT 204.600 128.800 205.000 129.200 ;
        RECT 204.600 127.200 204.900 128.800 ;
        RECT 204.600 126.800 205.000 127.200 ;
      LAYER via4 ;
        RECT 183.000 128.800 183.400 129.200 ;
      LAYER metal5 ;
        RECT 183.000 129.100 183.400 129.200 ;
        RECT 188.600 129.100 189.000 129.200 ;
        RECT 183.000 128.800 189.000 129.100 ;
    END
  END d_in[6]
  PIN d_in[7]
    PORT
      LAYER metal1 ;
        RECT 171.800 133.400 172.200 134.200 ;
        RECT 189.400 126.800 189.800 127.600 ;
      LAYER via1 ;
        RECT 171.800 133.800 172.200 134.200 ;
      LAYER metal2 ;
        RECT 171.800 133.800 172.200 134.200 ;
        RECT 171.800 131.200 172.100 133.800 ;
        RECT 171.800 130.800 172.200 131.200 ;
        RECT 188.600 130.800 189.000 131.200 ;
        RECT 188.600 127.100 188.900 130.800 ;
        RECT 189.400 127.100 189.800 127.200 ;
        RECT 188.600 126.800 189.800 127.100 ;
      LAYER metal3 ;
        RECT 171.800 131.100 172.200 131.200 ;
        RECT 188.600 131.100 189.000 131.200 ;
        RECT 207.800 131.100 208.200 131.200 ;
        RECT 171.800 130.800 208.200 131.100 ;
    END
  END d_in[7]
  PIN wr_en
    PORT
      LAYER metal1 ;
        RECT 193.400 175.400 193.800 176.200 ;
        RECT 190.600 156.800 191.000 157.200 ;
        RECT 190.700 156.200 191.000 156.800 ;
        RECT 190.700 155.900 191.400 156.200 ;
        RECT 191.000 155.800 191.400 155.900 ;
        RECT 193.400 154.800 193.800 155.200 ;
        RECT 193.400 154.400 193.700 154.800 ;
        RECT 193.200 154.100 193.700 154.400 ;
        RECT 193.200 154.000 193.600 154.100 ;
      LAYER via1 ;
        RECT 193.400 175.800 193.800 176.200 ;
      LAYER metal2 ;
        RECT 193.400 182.800 193.800 183.200 ;
        RECT 193.400 176.200 193.700 182.800 ;
        RECT 193.400 175.800 193.800 176.200 ;
        RECT 193.400 175.200 193.700 175.800 ;
        RECT 193.400 174.800 193.800 175.200 ;
        RECT 191.000 156.100 191.400 156.200 ;
        RECT 191.800 156.100 192.200 156.200 ;
        RECT 191.000 155.800 192.200 156.100 ;
        RECT 193.400 155.800 193.800 156.200 ;
        RECT 193.400 155.200 193.700 155.800 ;
        RECT 193.400 154.800 193.800 155.200 ;
      LAYER via2 ;
        RECT 191.800 155.800 192.200 156.200 ;
      LAYER metal3 ;
        RECT 193.400 175.800 193.800 176.200 ;
        RECT 193.400 175.200 193.700 175.800 ;
        RECT 193.400 174.800 193.800 175.200 ;
        RECT 191.800 156.100 192.200 156.200 ;
        RECT 193.400 156.100 193.800 156.200 ;
        RECT 191.800 155.800 193.800 156.100 ;
      LAYER via3 ;
        RECT 193.400 155.800 193.800 156.200 ;
      LAYER metal4 ;
        RECT 193.400 175.800 193.800 176.200 ;
        RECT 193.400 156.200 193.700 175.800 ;
        RECT 193.400 155.800 193.800 156.200 ;
    END
  END wr_en
  PIN rd_en
    PORT
      LAYER metal1 ;
        RECT 200.600 164.800 201.000 165.600 ;
        RECT 185.800 156.800 186.200 157.200 ;
        RECT 185.900 156.200 186.200 156.800 ;
        RECT 185.900 156.100 186.600 156.200 ;
        RECT 187.000 156.100 187.400 156.200 ;
        RECT 185.900 155.900 187.400 156.100 ;
        RECT 186.200 155.800 187.400 155.900 ;
        RECT 187.000 152.400 187.400 153.200 ;
        RECT 201.200 146.600 201.800 147.000 ;
        RECT 201.400 146.200 201.700 146.600 ;
        RECT 201.400 145.800 201.800 146.200 ;
        RECT 197.800 135.200 198.200 135.400 ;
        RECT 197.800 134.900 198.600 135.200 ;
        RECT 198.200 134.800 198.600 134.900 ;
      LAYER via1 ;
        RECT 187.000 155.800 187.400 156.200 ;
        RECT 187.000 152.800 187.400 153.200 ;
        RECT 201.400 146.600 201.800 147.000 ;
      LAYER metal2 ;
        RECT 195.800 182.800 196.200 183.200 ;
        RECT 195.800 171.200 196.100 182.800 ;
        RECT 195.800 170.800 196.200 171.200 ;
        RECT 200.600 170.800 201.000 171.200 ;
        RECT 200.600 165.200 200.900 170.800 ;
        RECT 200.600 164.800 201.000 165.200 ;
        RECT 187.000 155.800 187.400 156.200 ;
        RECT 187.000 153.200 187.300 155.800 ;
        RECT 200.600 153.200 200.900 164.800 ;
        RECT 187.000 153.100 187.400 153.200 ;
        RECT 187.800 153.100 188.200 153.200 ;
        RECT 187.000 152.800 188.200 153.100 ;
        RECT 200.600 152.800 201.000 153.200 ;
        RECT 200.600 151.100 200.900 152.800 ;
        RECT 200.600 150.800 201.700 151.100 ;
        RECT 200.600 135.200 200.900 150.800 ;
        RECT 201.400 147.000 201.700 150.800 ;
        RECT 201.400 146.600 201.800 147.000 ;
        RECT 198.200 135.100 198.600 135.200 ;
        RECT 199.000 135.100 199.400 135.200 ;
        RECT 198.200 134.800 199.400 135.100 ;
        RECT 200.600 134.800 201.000 135.200 ;
      LAYER via2 ;
        RECT 187.800 152.800 188.200 153.200 ;
        RECT 199.000 134.800 199.400 135.200 ;
      LAYER metal3 ;
        RECT 195.800 171.100 196.200 171.200 ;
        RECT 200.600 171.100 201.000 171.200 ;
        RECT 195.800 170.800 201.000 171.100 ;
        RECT 187.800 153.100 188.200 153.200 ;
        RECT 200.600 153.100 201.000 153.200 ;
        RECT 187.800 152.800 201.000 153.100 ;
        RECT 199.000 135.100 199.400 135.200 ;
        RECT 200.600 135.100 201.000 135.200 ;
        RECT 199.000 134.800 201.000 135.100 ;
    END
  END rd_en
  PIN full
    PORT
      LAYER metal1 ;
        RECT 199.800 177.100 200.200 179.900 ;
        RECT 199.800 176.800 200.900 177.100 ;
        RECT 199.800 175.900 200.200 176.800 ;
        RECT 199.900 174.800 200.200 175.900 ;
        RECT 200.600 176.200 200.900 176.800 ;
        RECT 200.600 175.800 201.000 176.200 ;
        RECT 199.800 171.100 200.200 174.800 ;
      LAYER metal2 ;
        RECT 200.600 176.800 201.000 177.200 ;
        RECT 200.600 176.200 200.900 176.800 ;
        RECT 200.600 175.800 201.000 176.200 ;
      LAYER metal3 ;
        RECT 200.600 177.100 201.000 177.200 ;
        RECT 207.800 177.100 208.200 177.200 ;
        RECT 200.600 176.800 208.200 177.100 ;
    END
  END full
  PIN empty
    PORT
      LAYER metal1 ;
        RECT 203.800 175.900 204.200 179.900 ;
        RECT 203.900 174.800 204.200 175.900 ;
        RECT 203.800 174.100 204.200 174.800 ;
        RECT 204.600 174.100 205.000 174.200 ;
        RECT 203.800 173.800 205.000 174.100 ;
        RECT 203.800 171.100 204.200 173.800 ;
      LAYER via1 ;
        RECT 204.600 173.800 205.000 174.200 ;
      LAYER metal2 ;
        RECT 204.600 174.800 205.000 175.200 ;
        RECT 204.600 174.200 204.900 174.800 ;
        RECT 204.600 173.800 205.000 174.200 ;
      LAYER metal3 ;
        RECT 204.600 175.100 205.000 175.200 ;
        RECT 207.800 175.100 208.200 175.200 ;
        RECT 204.600 174.800 208.200 175.100 ;
    END
  END empty
  PIN d_out[0]
    PORT
      LAYER metal1 ;
        RECT 3.000 155.900 3.400 159.900 ;
        RECT 3.000 154.800 3.300 155.900 ;
        RECT 3.000 151.100 3.400 154.800 ;
      LAYER via1 ;
        RECT 3.000 156.800 3.400 157.200 ;
      LAYER metal2 ;
        RECT 3.000 156.800 3.400 157.200 ;
        RECT 3.000 155.200 3.300 156.800 ;
        RECT 3.000 154.800 3.400 155.200 ;
      LAYER metal3 ;
        RECT -2.600 155.100 -2.200 155.200 ;
        RECT 3.000 155.100 3.400 155.200 ;
        RECT -2.600 154.800 3.400 155.100 ;
    END
  END d_out[0]
  PIN d_out[1]
    PORT
      LAYER metal1 ;
        RECT 0.600 155.900 1.000 159.900 ;
        RECT 0.600 154.800 0.900 155.900 ;
        RECT 0.600 151.100 1.000 154.800 ;
      LAYER via1 ;
        RECT 0.600 156.800 1.000 157.200 ;
      LAYER metal2 ;
        RECT 0.600 157.800 1.000 158.200 ;
        RECT 0.600 157.200 0.900 157.800 ;
        RECT 0.600 156.800 1.000 157.200 ;
      LAYER metal3 ;
        RECT 0.600 157.800 1.000 158.200 ;
        RECT -2.600 157.100 -2.200 157.200 ;
        RECT 0.600 157.100 0.900 157.800 ;
        RECT -2.600 156.800 0.900 157.100 ;
    END
  END d_out[1]
  PIN d_out[2]
    PORT
      LAYER metal1 ;
        RECT 40.600 175.900 41.000 179.900 ;
        RECT 40.600 174.800 40.900 175.900 ;
        RECT 40.600 171.100 41.000 174.800 ;
      LAYER via1 ;
        RECT 40.600 171.800 41.000 172.200 ;
      LAYER metal2 ;
        RECT 40.600 172.800 41.000 173.200 ;
        RECT 40.600 172.200 40.900 172.800 ;
        RECT 40.600 171.800 41.000 172.200 ;
      LAYER metal3 ;
        RECT 40.600 172.800 41.000 173.200 ;
        RECT -2.600 172.100 -2.200 172.200 ;
        RECT 40.600 172.100 40.900 172.800 ;
        RECT -2.600 171.800 40.900 172.100 ;
    END
  END d_out[2]
  PIN d_out[3]
    PORT
      LAYER metal1 ;
        RECT 15.000 175.900 15.400 179.900 ;
        RECT 15.000 174.800 15.300 175.900 ;
        RECT 15.000 171.100 15.400 174.800 ;
      LAYER via1 ;
        RECT 15.000 173.800 15.400 174.200 ;
      LAYER metal2 ;
        RECT 15.000 174.800 15.400 175.200 ;
        RECT 15.000 174.200 15.300 174.800 ;
        RECT 15.000 173.800 15.400 174.200 ;
      LAYER metal3 ;
        RECT 15.000 175.100 15.400 175.200 ;
        RECT 1.400 174.800 15.400 175.100 ;
        RECT -2.600 174.100 -2.200 174.200 ;
        RECT 1.400 174.100 1.700 174.800 ;
        RECT -2.600 173.800 1.700 174.100 ;
    END
  END d_out[3]
  PIN d_out[4]
    PORT
      LAYER metal1 ;
        RECT 12.600 175.900 13.000 179.900 ;
        RECT 12.600 174.800 12.900 175.900 ;
        RECT 12.600 171.100 13.000 174.800 ;
      LAYER via1 ;
        RECT 12.600 173.800 13.000 174.200 ;
      LAYER metal2 ;
        RECT 12.600 175.800 13.000 176.200 ;
        RECT 12.600 174.200 12.900 175.800 ;
        RECT 12.600 173.800 13.000 174.200 ;
      LAYER metal3 ;
        RECT -2.600 176.100 -2.200 176.200 ;
        RECT 12.600 176.100 13.000 176.200 ;
        RECT -2.600 175.800 13.000 176.100 ;
    END
  END d_out[4]
  PIN d_out[5]
    PORT
      LAYER metal1 ;
        RECT 17.400 175.900 17.800 179.900 ;
        RECT 17.400 174.800 17.700 175.900 ;
        RECT 17.400 171.100 17.800 174.800 ;
      LAYER via1 ;
        RECT 17.400 178.800 17.800 179.200 ;
      LAYER metal2 ;
        RECT 17.400 179.800 17.800 180.200 ;
        RECT 17.400 179.200 17.700 179.800 ;
        RECT 17.400 178.800 17.800 179.200 ;
      LAYER metal3 ;
        RECT 0.600 180.100 1.000 180.200 ;
        RECT 17.400 180.100 17.800 180.200 ;
        RECT 0.600 179.800 17.800 180.100 ;
        RECT -2.600 178.100 -2.200 178.200 ;
        RECT 0.600 178.100 1.000 178.200 ;
        RECT -2.600 177.800 1.000 178.100 ;
      LAYER via3 ;
        RECT 0.600 177.800 1.000 178.200 ;
      LAYER metal4 ;
        RECT 0.600 179.800 1.000 180.200 ;
        RECT 0.600 178.200 0.900 179.800 ;
        RECT 0.600 177.800 1.000 178.200 ;
    END
  END d_out[5]
  PIN d_out[6]
    PORT
      LAYER metal1 ;
        RECT 0.600 175.900 1.000 179.900 ;
        RECT 0.600 174.800 0.900 175.900 ;
        RECT 0.600 171.100 1.000 174.800 ;
      LAYER via1 ;
        RECT 0.600 178.800 1.000 179.200 ;
      LAYER metal2 ;
        RECT 0.600 179.100 1.000 179.200 ;
        RECT 1.400 179.100 1.800 179.200 ;
        RECT 0.600 178.800 1.800 179.100 ;
      LAYER via2 ;
        RECT 1.400 178.800 1.800 179.200 ;
      LAYER metal3 ;
        RECT -2.600 179.800 -2.200 180.200 ;
        RECT -2.600 179.100 -2.300 179.800 ;
        RECT 1.400 179.100 1.800 179.200 ;
        RECT -2.600 178.800 1.800 179.100 ;
    END
  END d_out[6]
  PIN d_out[7]
    PORT
      LAYER metal1 ;
        RECT 3.000 175.900 3.400 179.900 ;
        RECT 3.000 174.800 3.300 175.900 ;
        RECT 3.000 171.100 3.400 174.800 ;
      LAYER via1 ;
        RECT 3.000 178.800 3.400 179.200 ;
      LAYER metal2 ;
        RECT 3.000 178.800 3.400 179.200 ;
        RECT 3.000 178.200 3.300 178.800 ;
        RECT 3.000 177.800 3.400 178.200 ;
      LAYER metal3 ;
        RECT -2.600 181.800 -2.200 182.200 ;
        RECT 2.200 179.100 2.600 179.200 ;
        RECT 2.200 178.800 3.300 179.100 ;
        RECT 3.000 178.200 3.300 178.800 ;
        RECT 3.000 177.800 3.400 178.200 ;
      LAYER metal4 ;
        RECT -2.600 182.100 -2.200 182.200 ;
        RECT -1.800 182.100 -1.400 182.200 ;
        RECT -2.600 181.800 -1.400 182.100 ;
        RECT 2.200 179.800 2.600 180.200 ;
        RECT 2.200 179.200 2.500 179.800 ;
        RECT 2.200 178.800 2.600 179.200 ;
      LAYER via4 ;
        RECT -1.800 181.800 -1.400 182.200 ;
      LAYER metal5 ;
        RECT -1.800 182.100 -1.400 182.200 ;
        RECT -2.600 181.800 -1.400 182.100 ;
        RECT -2.600 180.100 -2.300 181.800 ;
        RECT 2.200 180.100 2.600 180.200 ;
        RECT -2.600 179.800 2.600 180.100 ;
    END
  END d_out[7]
  PIN fifo_counter[0]
    PORT
      LAYER metal1 ;
        RECT 199.800 26.200 200.200 29.900 ;
        RECT 199.800 25.100 200.100 26.200 ;
        RECT 199.800 21.100 200.200 25.100 ;
      LAYER via1 ;
        RECT 199.800 21.800 200.200 22.200 ;
      LAYER metal2 ;
        RECT 199.800 21.800 200.200 22.200 ;
        RECT 199.800 20.200 200.100 21.800 ;
        RECT 199.800 19.800 200.200 20.200 ;
        RECT 199.000 0.800 199.400 1.200 ;
        RECT 199.000 -1.800 199.300 0.800 ;
        RECT 199.000 -2.200 199.400 -1.800 ;
      LAYER metal3 ;
        RECT 199.000 20.100 199.400 20.200 ;
        RECT 199.800 20.100 200.200 20.200 ;
        RECT 199.000 19.800 200.200 20.100 ;
        RECT 199.000 1.100 199.400 1.200 ;
        RECT 199.800 1.100 200.200 1.200 ;
        RECT 199.000 0.800 200.200 1.100 ;
      LAYER via3 ;
        RECT 199.800 0.800 200.200 1.200 ;
      LAYER metal4 ;
        RECT 199.000 19.800 199.400 20.200 ;
        RECT 199.000 1.100 199.300 19.800 ;
        RECT 199.800 1.100 200.200 1.200 ;
        RECT 199.000 0.800 200.200 1.100 ;
    END
  END fifo_counter[0]
  PIN fifo_counter[1]
    PORT
      LAYER metal1 ;
        RECT 203.000 146.200 203.400 149.900 ;
        RECT 203.000 145.100 203.300 146.200 ;
        RECT 203.000 141.100 203.400 145.100 ;
      LAYER via1 ;
        RECT 203.000 141.800 203.400 142.200 ;
      LAYER metal2 ;
        RECT 203.000 141.800 203.400 142.200 ;
        RECT 203.000 137.100 203.300 141.800 ;
        RECT 203.800 137.100 204.200 137.200 ;
        RECT 203.000 136.800 204.200 137.100 ;
        RECT 201.400 0.800 201.800 1.200 ;
        RECT 201.400 -1.800 201.700 0.800 ;
        RECT 201.400 -2.200 201.800 -1.800 ;
      LAYER via2 ;
        RECT 203.800 136.800 204.200 137.200 ;
      LAYER metal3 ;
        RECT 203.000 137.100 203.400 137.200 ;
        RECT 203.800 137.100 204.200 137.200 ;
        RECT 203.000 136.800 204.200 137.100 ;
        RECT 201.400 1.100 201.800 1.200 ;
        RECT 203.000 1.100 203.400 1.200 ;
        RECT 201.400 0.800 203.400 1.100 ;
      LAYER via3 ;
        RECT 203.000 0.800 203.400 1.200 ;
      LAYER metal4 ;
        RECT 203.000 136.800 203.400 137.200 ;
        RECT 203.000 1.200 203.300 136.800 ;
        RECT 203.000 0.800 203.400 1.200 ;
    END
  END fifo_counter[1]
  PIN fifo_counter[2]
    PORT
      LAYER metal1 ;
        RECT 203.000 15.900 203.400 19.900 ;
        RECT 203.100 14.800 203.400 15.900 ;
        RECT 203.000 12.100 203.400 14.800 ;
        RECT 203.800 12.100 204.200 12.200 ;
        RECT 203.000 11.800 204.200 12.100 ;
        RECT 203.000 11.100 203.400 11.800 ;
      LAYER via1 ;
        RECT 203.800 11.800 204.200 12.200 ;
      LAYER metal2 ;
        RECT 203.800 11.800 204.200 12.200 ;
        RECT 203.000 -1.900 203.400 -1.800 ;
        RECT 203.800 -1.900 204.100 11.800 ;
        RECT 203.000 -2.200 204.100 -1.900 ;
    END
  END fifo_counter[2]
  PIN fifo_counter[3]
    PORT
      LAYER metal1 ;
        RECT 199.000 15.900 199.400 19.900 ;
        RECT 199.100 14.800 199.400 15.900 ;
        RECT 199.000 11.100 199.400 14.800 ;
      LAYER via1 ;
        RECT 199.000 11.800 199.400 12.200 ;
      LAYER metal2 ;
        RECT 199.000 11.800 199.400 12.200 ;
        RECT 199.000 10.200 199.300 11.800 ;
        RECT 199.000 9.800 199.400 10.200 ;
        RECT 201.400 9.800 201.800 10.200 ;
        RECT 201.400 2.100 201.700 9.800 ;
        RECT 201.400 1.800 202.500 2.100 ;
        RECT 202.200 -2.900 202.500 1.800 ;
        RECT 204.600 -2.200 205.000 -1.800 ;
        RECT 204.600 -2.900 204.900 -2.200 ;
        RECT 202.200 -3.200 204.900 -2.900 ;
      LAYER metal3 ;
        RECT 199.000 10.100 199.400 10.200 ;
        RECT 201.400 10.100 201.800 10.200 ;
        RECT 199.000 9.800 201.800 10.100 ;
    END
  END fifo_counter[3]
  PIN fifo_counter[4]
    PORT
      LAYER metal1 ;
        RECT 203.800 26.200 204.200 29.900 ;
        RECT 203.900 25.100 204.200 26.200 ;
        RECT 203.800 22.100 204.200 25.100 ;
        RECT 204.600 22.100 205.000 22.200 ;
        RECT 203.800 21.800 205.000 22.100 ;
        RECT 203.800 21.100 204.200 21.800 ;
      LAYER via1 ;
        RECT 204.600 21.800 205.000 22.200 ;
      LAYER metal2 ;
        RECT 204.600 21.800 205.000 22.200 ;
        RECT 204.600 -0.900 204.900 21.800 ;
        RECT 204.600 -1.200 205.700 -0.900 ;
        RECT 205.400 -1.900 205.700 -1.200 ;
        RECT 206.200 -1.900 206.600 -1.800 ;
        RECT 205.400 -2.200 206.600 -1.900 ;
    END
  END fifo_counter[4]
  OBS
      LAYER metal1 ;
        RECT 2.200 176.200 2.600 179.900 ;
        RECT 4.600 176.200 5.000 179.900 ;
        RECT 1.500 175.900 2.600 176.200 ;
        RECT 3.900 175.900 5.000 176.200 ;
        RECT 1.500 175.600 1.800 175.900 ;
        RECT 3.900 175.600 4.200 175.900 ;
        RECT 1.200 175.200 1.800 175.600 ;
        RECT 3.600 175.200 4.200 175.600 ;
        RECT 6.200 175.600 6.600 179.900 ;
        RECT 7.800 175.600 8.200 179.900 ;
        RECT 9.400 175.600 9.800 179.900 ;
        RECT 11.000 175.600 11.400 179.900 ;
        RECT 14.200 176.200 14.600 179.900 ;
        RECT 16.600 176.200 17.000 179.900 ;
        RECT 19.000 176.200 19.400 179.900 ;
        RECT 13.500 175.900 14.600 176.200 ;
        RECT 15.900 175.900 17.000 176.200 ;
        RECT 18.300 175.900 19.400 176.200 ;
        RECT 20.600 176.000 21.000 179.900 ;
        RECT 22.200 177.600 22.600 179.900 ;
        RECT 13.500 175.600 13.800 175.900 ;
        RECT 15.900 175.600 16.200 175.900 ;
        RECT 18.300 175.600 18.600 175.900 ;
        RECT 6.200 175.200 7.100 175.600 ;
        RECT 7.800 175.200 8.900 175.600 ;
        RECT 9.400 175.200 10.500 175.600 ;
        RECT 11.000 175.200 12.200 175.600 ;
        RECT 13.200 175.200 13.800 175.600 ;
        RECT 15.600 175.200 16.200 175.600 ;
        RECT 18.000 175.200 18.600 175.600 ;
        RECT 20.500 175.600 21.000 176.000 ;
        RECT 21.300 177.300 22.600 177.600 ;
        RECT 21.300 176.500 21.600 177.300 ;
        RECT 23.800 177.200 24.200 179.900 ;
        RECT 25.400 178.500 25.800 179.900 ;
        RECT 26.200 178.500 26.600 179.900 ;
        RECT 27.000 178.500 27.400 179.900 ;
        RECT 24.500 177.200 26.600 177.600 ;
        RECT 22.900 176.800 24.200 177.200 ;
        RECT 27.800 176.800 28.200 179.900 ;
        RECT 29.400 177.500 29.800 179.900 ;
        RECT 31.000 177.500 31.400 179.900 ;
        RECT 31.800 178.500 32.200 179.900 ;
        RECT 32.600 178.500 33.000 179.900 ;
        RECT 34.200 177.600 34.600 179.900 ;
        RECT 35.800 178.200 36.200 179.900 ;
        RECT 35.800 177.900 36.300 178.200 ;
        RECT 36.000 177.600 36.300 177.900 ;
        RECT 33.600 177.200 35.700 177.600 ;
        RECT 36.000 177.300 37.000 177.600 ;
        RECT 29.400 176.800 30.700 177.200 ;
        RECT 31.000 176.900 33.900 177.200 ;
        RECT 35.400 177.000 35.700 177.200 ;
        RECT 25.400 176.500 25.800 176.600 ;
        RECT 21.300 176.200 25.800 176.500 ;
        RECT 27.000 176.500 27.400 176.600 ;
        RECT 31.000 176.500 31.300 176.900 ;
        RECT 34.200 176.600 34.900 176.900 ;
        RECT 35.400 176.600 36.200 177.000 ;
        RECT 27.000 176.200 31.300 176.500 ;
        RECT 31.800 176.500 34.900 176.600 ;
        RECT 31.800 176.300 34.500 176.500 ;
        RECT 31.800 176.200 32.200 176.300 ;
        RECT 1.500 173.700 1.800 175.200 ;
        RECT 2.200 174.400 2.600 175.200 ;
        RECT 3.900 173.700 4.200 175.200 ;
        RECT 4.600 174.400 5.000 175.200 ;
        RECT 6.700 174.500 7.100 175.200 ;
        RECT 8.500 174.500 8.900 175.200 ;
        RECT 10.100 174.500 10.500 175.200 ;
        RECT 6.700 174.100 8.000 174.500 ;
        RECT 8.500 174.100 9.700 174.500 ;
        RECT 10.100 174.100 11.400 174.500 ;
        RECT 6.700 173.800 7.100 174.100 ;
        RECT 8.500 173.800 8.900 174.100 ;
        RECT 10.100 173.800 10.500 174.100 ;
        RECT 11.800 173.800 12.200 175.200 ;
        RECT 1.500 173.400 2.600 173.700 ;
        RECT 3.900 173.400 5.000 173.700 ;
        RECT 2.200 171.100 2.600 173.400 ;
        RECT 4.600 171.100 5.000 173.400 ;
        RECT 6.200 173.400 7.100 173.800 ;
        RECT 7.800 173.400 8.900 173.800 ;
        RECT 9.400 173.400 10.500 173.800 ;
        RECT 11.000 173.400 12.200 173.800 ;
        RECT 13.500 173.700 13.800 175.200 ;
        RECT 14.200 174.400 14.600 175.200 ;
        RECT 15.900 173.700 16.200 175.200 ;
        RECT 16.600 174.400 17.000 175.200 ;
        RECT 18.300 173.700 18.600 175.200 ;
        RECT 19.000 175.100 19.400 175.200 ;
        RECT 20.500 175.100 20.900 175.600 ;
        RECT 21.300 175.300 21.600 176.200 ;
        RECT 19.000 174.800 20.900 175.100 ;
        RECT 19.000 174.400 19.400 174.800 ;
        RECT 13.500 173.400 14.600 173.700 ;
        RECT 15.900 173.400 17.000 173.700 ;
        RECT 18.300 173.400 19.400 173.700 ;
        RECT 6.200 171.100 6.600 173.400 ;
        RECT 7.800 171.100 8.200 173.400 ;
        RECT 9.400 171.100 9.800 173.400 ;
        RECT 11.000 171.100 11.400 173.400 ;
        RECT 14.200 171.100 14.600 173.400 ;
        RECT 16.600 171.100 17.000 173.400 ;
        RECT 19.000 171.100 19.400 173.400 ;
        RECT 20.500 173.400 20.900 174.800 ;
        RECT 21.200 175.000 21.600 175.300 ;
        RECT 24.600 175.000 36.300 175.300 ;
        RECT 21.200 174.000 21.500 175.000 ;
        RECT 24.600 174.700 25.000 175.000 ;
        RECT 33.400 174.800 33.800 175.000 ;
        RECT 35.000 174.800 35.400 175.000 ;
        RECT 35.900 174.900 36.300 175.000 ;
        RECT 21.800 174.300 23.700 174.700 ;
        RECT 21.200 173.700 21.800 174.000 ;
        RECT 20.500 173.000 21.000 173.400 ;
        RECT 20.600 171.100 21.000 173.000 ;
        RECT 21.400 171.100 21.800 173.700 ;
        RECT 23.300 173.700 23.700 174.300 ;
        RECT 23.300 173.400 24.200 173.700 ;
        RECT 23.800 173.100 24.200 173.400 ;
        RECT 26.200 173.200 26.600 174.600 ;
        RECT 27.800 174.300 29.400 174.700 ;
        RECT 31.300 174.300 32.300 174.700 ;
        RECT 36.600 174.500 37.000 177.300 ;
        RECT 38.200 176.400 38.600 179.900 ;
        RECT 38.100 175.900 38.600 176.400 ;
        RECT 39.800 176.200 40.200 179.900 ;
        RECT 42.200 176.200 42.600 179.900 ;
        RECT 38.900 175.900 40.200 176.200 ;
        RECT 41.500 175.900 42.600 176.200 ;
        RECT 45.400 176.000 45.800 179.900 ;
        RECT 47.000 177.600 47.400 179.900 ;
        RECT 27.600 173.900 28.000 174.000 ;
        RECT 27.600 173.600 29.800 173.900 ;
        RECT 29.400 173.500 29.800 173.600 ;
        RECT 30.200 173.400 30.600 174.200 ;
        RECT 23.800 172.700 25.000 173.100 ;
        RECT 26.200 172.800 26.700 173.200 ;
        RECT 28.200 172.800 29.000 173.200 ;
        RECT 29.400 173.100 29.800 173.200 ;
        RECT 31.300 173.100 31.700 174.300 ;
        RECT 32.600 174.100 37.000 174.500 ;
        RECT 34.300 173.400 35.800 173.800 ;
        RECT 34.300 173.100 34.700 173.400 ;
        RECT 29.400 172.800 31.700 173.100 ;
        RECT 24.600 171.100 25.000 172.700 ;
        RECT 33.400 172.700 34.700 173.100 ;
        RECT 25.400 171.100 25.800 172.500 ;
        RECT 26.200 171.100 26.600 172.500 ;
        RECT 27.000 171.100 27.400 172.500 ;
        RECT 27.800 171.100 28.200 172.500 ;
        RECT 29.400 171.100 29.800 172.500 ;
        RECT 31.000 171.100 31.400 172.500 ;
        RECT 31.800 171.100 32.200 172.500 ;
        RECT 32.600 171.100 33.000 172.500 ;
        RECT 33.400 171.100 33.800 172.700 ;
        RECT 36.600 171.100 37.000 174.100 ;
        RECT 37.400 174.800 37.800 175.200 ;
        RECT 37.400 174.100 37.700 174.800 ;
        RECT 38.100 174.200 38.400 175.900 ;
        RECT 38.900 174.900 39.200 175.900 ;
        RECT 41.500 175.600 41.800 175.900 ;
        RECT 41.200 175.200 41.800 175.600 ;
        RECT 45.300 175.600 45.800 176.000 ;
        RECT 46.100 177.300 47.400 177.600 ;
        RECT 46.100 176.500 46.400 177.300 ;
        RECT 48.600 177.200 49.000 179.900 ;
        RECT 50.200 178.500 50.600 179.900 ;
        RECT 51.000 178.500 51.400 179.900 ;
        RECT 51.800 178.500 52.200 179.900 ;
        RECT 49.300 177.200 51.400 177.600 ;
        RECT 47.700 176.800 49.000 177.200 ;
        RECT 52.600 176.800 53.000 179.900 ;
        RECT 54.200 177.500 54.600 179.900 ;
        RECT 55.800 177.500 56.200 179.900 ;
        RECT 56.600 178.500 57.000 179.900 ;
        RECT 57.400 178.500 57.800 179.900 ;
        RECT 59.000 177.600 59.400 179.900 ;
        RECT 60.600 178.200 61.000 179.900 ;
        RECT 60.600 177.900 61.100 178.200 ;
        RECT 60.800 177.600 61.100 177.900 ;
        RECT 58.400 177.200 60.500 177.600 ;
        RECT 60.800 177.300 61.800 177.600 ;
        RECT 54.200 176.800 55.500 177.200 ;
        RECT 55.800 176.900 58.700 177.200 ;
        RECT 60.200 177.000 60.500 177.200 ;
        RECT 50.200 176.500 50.600 176.600 ;
        RECT 46.100 176.200 50.600 176.500 ;
        RECT 51.800 176.500 52.200 176.600 ;
        RECT 55.800 176.500 56.100 176.900 ;
        RECT 59.000 176.600 59.700 176.900 ;
        RECT 60.200 176.600 61.000 177.000 ;
        RECT 51.800 176.200 56.100 176.500 ;
        RECT 56.600 176.500 59.700 176.600 ;
        RECT 56.600 176.300 59.300 176.500 ;
        RECT 56.600 176.200 57.000 176.300 ;
        RECT 38.700 174.500 39.200 174.900 ;
        RECT 38.100 174.100 38.600 174.200 ;
        RECT 37.400 173.800 38.600 174.100 ;
        RECT 38.100 173.100 38.400 173.800 ;
        RECT 38.900 173.700 39.200 174.500 ;
        RECT 39.700 174.800 40.200 175.200 ;
        RECT 39.700 174.400 40.100 174.800 ;
        RECT 41.500 173.700 41.800 175.200 ;
        RECT 42.200 175.100 42.600 175.200 ;
        RECT 45.300 175.100 45.700 175.600 ;
        RECT 46.100 175.300 46.400 176.200 ;
        RECT 42.200 174.800 45.700 175.100 ;
        RECT 42.200 174.400 42.600 174.800 ;
        RECT 38.900 173.400 40.200 173.700 ;
        RECT 41.500 173.400 42.600 173.700 ;
        RECT 38.100 172.800 38.600 173.100 ;
        RECT 38.200 171.100 38.600 172.800 ;
        RECT 39.800 171.100 40.200 173.400 ;
        RECT 42.200 171.100 42.600 173.400 ;
        RECT 45.300 173.400 45.700 174.800 ;
        RECT 46.000 175.000 46.400 175.300 ;
        RECT 49.400 175.000 61.100 175.300 ;
        RECT 46.000 174.000 46.300 175.000 ;
        RECT 49.400 174.700 49.800 175.000 ;
        RECT 58.200 174.800 58.600 175.000 ;
        RECT 60.700 174.900 61.100 175.000 ;
        RECT 46.600 174.300 48.500 174.700 ;
        RECT 46.000 173.700 46.600 174.000 ;
        RECT 45.300 173.000 45.800 173.400 ;
        RECT 45.400 171.100 45.800 173.000 ;
        RECT 46.200 171.100 46.600 173.700 ;
        RECT 48.100 173.700 48.500 174.300 ;
        RECT 48.100 173.400 49.000 173.700 ;
        RECT 48.600 173.100 49.000 173.400 ;
        RECT 51.000 173.200 51.400 174.600 ;
        RECT 52.600 174.300 54.200 174.700 ;
        RECT 56.100 174.300 57.100 174.700 ;
        RECT 61.400 174.500 61.800 177.300 ;
        RECT 52.400 173.900 52.800 174.000 ;
        RECT 52.400 173.600 54.600 173.900 ;
        RECT 54.200 173.500 54.600 173.600 ;
        RECT 55.000 173.400 55.400 174.200 ;
        RECT 48.600 172.700 49.800 173.100 ;
        RECT 51.000 172.800 51.500 173.200 ;
        RECT 53.000 172.800 53.800 173.200 ;
        RECT 54.200 173.100 54.600 173.200 ;
        RECT 56.100 173.100 56.500 174.300 ;
        RECT 57.400 174.100 61.800 174.500 ;
        RECT 59.100 173.400 60.600 173.800 ;
        RECT 59.100 173.100 59.500 173.400 ;
        RECT 54.200 172.800 56.500 173.100 ;
        RECT 49.400 171.100 49.800 172.700 ;
        RECT 58.200 172.700 59.500 173.100 ;
        RECT 50.200 171.100 50.600 172.500 ;
        RECT 51.000 171.100 51.400 172.500 ;
        RECT 51.800 171.100 52.200 172.500 ;
        RECT 52.600 171.100 53.000 172.500 ;
        RECT 54.200 171.100 54.600 172.500 ;
        RECT 55.800 171.100 56.200 172.500 ;
        RECT 56.600 171.100 57.000 172.500 ;
        RECT 57.400 171.100 57.800 172.500 ;
        RECT 58.200 171.100 58.600 172.700 ;
        RECT 61.400 171.100 61.800 174.100 ;
        RECT 62.200 175.600 62.600 179.900 ;
        RECT 64.300 177.900 64.900 179.900 ;
        RECT 66.600 177.900 67.000 179.900 ;
        RECT 68.800 178.200 69.200 179.900 ;
        RECT 68.800 177.900 69.800 178.200 ;
        RECT 64.600 177.500 65.000 177.900 ;
        RECT 66.700 177.600 67.000 177.900 ;
        RECT 66.300 177.300 68.100 177.600 ;
        RECT 69.400 177.500 69.800 177.900 ;
        RECT 66.300 177.200 66.700 177.300 ;
        RECT 67.700 177.200 68.100 177.300 ;
        RECT 64.200 176.600 64.900 177.000 ;
        RECT 64.600 176.100 64.900 176.600 ;
        RECT 65.700 176.500 66.800 176.800 ;
        RECT 65.700 176.400 66.100 176.500 ;
        RECT 64.600 175.800 65.800 176.100 ;
        RECT 62.200 175.300 64.300 175.600 ;
        RECT 62.200 173.600 62.600 175.300 ;
        RECT 63.900 175.200 64.300 175.300 ;
        RECT 63.100 174.900 63.500 175.000 ;
        RECT 63.100 174.600 65.000 174.900 ;
        RECT 64.600 174.500 65.000 174.600 ;
        RECT 65.500 174.200 65.800 175.800 ;
        RECT 66.500 175.900 66.800 176.500 ;
        RECT 67.100 176.500 67.500 176.600 ;
        RECT 69.400 176.500 69.800 176.600 ;
        RECT 67.100 176.200 69.800 176.500 ;
        RECT 66.500 175.700 68.900 175.900 ;
        RECT 71.000 175.700 71.400 179.900 ;
        RECT 66.500 175.600 71.400 175.700 ;
        RECT 68.500 175.500 71.400 175.600 ;
        RECT 68.600 175.400 71.400 175.500 ;
        RECT 71.800 175.600 72.200 179.900 ;
        RECT 73.900 177.900 74.500 179.900 ;
        RECT 76.200 177.900 76.600 179.900 ;
        RECT 78.400 178.200 78.800 179.900 ;
        RECT 78.400 177.900 79.400 178.200 ;
        RECT 74.200 177.500 74.600 177.900 ;
        RECT 76.300 177.600 76.600 177.900 ;
        RECT 75.900 177.300 77.700 177.600 ;
        RECT 79.000 177.500 79.400 177.900 ;
        RECT 75.900 177.200 76.300 177.300 ;
        RECT 77.300 177.200 77.700 177.300 ;
        RECT 73.800 176.600 74.500 177.000 ;
        RECT 74.200 176.100 74.500 176.600 ;
        RECT 75.300 176.500 76.400 176.800 ;
        RECT 75.300 176.400 75.700 176.500 ;
        RECT 74.200 175.800 75.400 176.100 ;
        RECT 71.800 175.300 73.900 175.600 ;
        RECT 67.800 175.100 68.200 175.200 ;
        RECT 67.800 174.800 70.300 175.100 ;
        RECT 69.900 174.700 70.300 174.800 ;
        RECT 69.100 174.200 69.500 174.300 ;
        RECT 65.500 173.900 71.000 174.200 ;
        RECT 65.700 173.800 66.600 173.900 ;
        RECT 62.200 173.300 64.100 173.600 ;
        RECT 62.200 171.100 62.600 173.300 ;
        RECT 63.700 173.200 64.100 173.300 ;
        RECT 68.600 172.800 68.900 173.900 ;
        RECT 70.200 173.800 71.000 173.900 ;
        RECT 71.800 173.600 72.200 175.300 ;
        RECT 73.500 175.200 73.900 175.300 ;
        RECT 72.700 174.900 73.100 175.000 ;
        RECT 72.700 174.600 74.600 174.900 ;
        RECT 74.200 174.500 74.600 174.600 ;
        RECT 75.100 174.200 75.400 175.800 ;
        RECT 76.100 175.900 76.400 176.500 ;
        RECT 76.700 176.500 77.100 176.600 ;
        RECT 79.000 176.500 79.400 176.600 ;
        RECT 76.700 176.200 79.400 176.500 ;
        RECT 76.100 175.700 78.500 175.900 ;
        RECT 80.600 175.700 81.000 179.900 ;
        RECT 76.100 175.600 81.000 175.700 ;
        RECT 78.100 175.500 81.000 175.600 ;
        RECT 78.200 175.400 81.000 175.500 ;
        RECT 82.200 175.600 82.600 179.900 ;
        RECT 83.800 175.600 84.200 179.900 ;
        RECT 86.200 175.600 86.600 179.900 ;
        RECT 87.800 175.600 88.200 179.900 ;
        RECT 89.400 175.600 89.800 179.900 ;
        RECT 91.000 175.600 91.400 179.900 ;
        RECT 93.400 178.200 93.800 179.900 ;
        RECT 93.300 177.900 93.800 178.200 ;
        RECT 93.300 177.600 93.600 177.900 ;
        RECT 95.000 177.600 95.400 179.900 ;
        RECT 96.600 178.500 97.000 179.900 ;
        RECT 97.400 178.500 97.800 179.900 ;
        RECT 82.200 175.200 84.200 175.600 ;
        RECT 77.400 175.100 77.800 175.200 ;
        RECT 77.400 174.800 79.900 175.100 ;
        RECT 79.500 174.700 79.900 174.800 ;
        RECT 78.700 174.200 79.100 174.300 ;
        RECT 75.000 173.900 80.600 174.200 ;
        RECT 75.000 173.800 75.700 173.900 ;
        RECT 67.700 172.700 68.100 172.800 ;
        RECT 64.600 172.100 65.000 172.500 ;
        RECT 66.700 172.400 68.100 172.700 ;
        RECT 68.600 172.400 69.000 172.800 ;
        RECT 66.700 172.100 67.000 172.400 ;
        RECT 69.400 172.100 69.800 172.500 ;
        RECT 64.300 171.800 65.000 172.100 ;
        RECT 64.300 171.100 64.900 171.800 ;
        RECT 66.600 171.100 67.000 172.100 ;
        RECT 68.800 171.800 69.800 172.100 ;
        RECT 68.800 171.100 69.200 171.800 ;
        RECT 71.000 171.100 71.400 173.500 ;
        RECT 71.800 173.300 73.700 173.600 ;
        RECT 71.800 171.100 72.200 173.300 ;
        RECT 73.300 173.200 73.700 173.300 ;
        RECT 78.200 172.800 78.500 173.900 ;
        RECT 79.800 173.800 80.600 173.900 ;
        RECT 83.800 173.800 84.200 175.200 ;
        RECT 85.400 175.200 86.600 175.600 ;
        RECT 87.100 175.200 88.200 175.600 ;
        RECT 88.700 175.200 89.800 175.600 ;
        RECT 90.500 175.200 91.400 175.600 ;
        RECT 92.600 177.300 93.600 177.600 ;
        RECT 84.600 174.100 85.000 174.200 ;
        RECT 85.400 174.100 85.800 175.200 ;
        RECT 87.100 174.500 87.500 175.200 ;
        RECT 88.700 174.500 89.100 175.200 ;
        RECT 90.500 174.500 90.900 175.200 ;
        RECT 86.200 174.100 87.500 174.500 ;
        RECT 87.900 174.100 89.100 174.500 ;
        RECT 89.600 174.100 90.900 174.500 ;
        RECT 84.600 173.800 85.800 174.100 ;
        RECT 87.100 173.800 87.500 174.100 ;
        RECT 88.700 173.800 89.100 174.100 ;
        RECT 90.500 173.800 90.900 174.100 ;
        RECT 92.600 174.500 93.000 177.300 ;
        RECT 93.900 177.200 96.000 177.600 ;
        RECT 98.200 177.500 98.600 179.900 ;
        RECT 99.800 177.500 100.200 179.900 ;
        RECT 93.900 177.000 94.200 177.200 ;
        RECT 93.400 176.600 94.200 177.000 ;
        RECT 95.700 176.900 98.600 177.200 ;
        RECT 94.700 176.600 95.400 176.900 ;
        RECT 94.700 176.500 97.800 176.600 ;
        RECT 95.100 176.300 97.800 176.500 ;
        RECT 97.400 176.200 97.800 176.300 ;
        RECT 98.300 176.500 98.600 176.900 ;
        RECT 98.900 176.800 100.200 177.200 ;
        RECT 101.400 176.800 101.800 179.900 ;
        RECT 102.200 178.500 102.600 179.900 ;
        RECT 103.000 178.500 103.400 179.900 ;
        RECT 103.800 178.500 104.200 179.900 ;
        RECT 103.000 177.200 105.100 177.600 ;
        RECT 105.400 177.200 105.800 179.900 ;
        RECT 107.000 177.600 107.400 179.900 ;
        RECT 107.000 177.300 108.300 177.600 ;
        RECT 105.400 176.800 106.700 177.200 ;
        RECT 102.200 176.500 102.600 176.600 ;
        RECT 98.300 176.200 102.600 176.500 ;
        RECT 103.800 176.500 104.200 176.600 ;
        RECT 108.000 176.500 108.300 177.300 ;
        RECT 103.800 176.200 108.300 176.500 ;
        RECT 108.000 175.300 108.300 176.200 ;
        RECT 108.600 176.000 109.000 179.900 ;
        RECT 111.800 176.200 112.200 179.900 ;
        RECT 113.400 176.400 113.800 179.900 ;
        RECT 108.600 175.600 109.100 176.000 ;
        RECT 111.800 175.900 113.100 176.200 ;
        RECT 113.400 175.900 113.900 176.400 ;
        RECT 93.300 175.000 105.000 175.300 ;
        RECT 108.000 175.000 108.400 175.300 ;
        RECT 93.300 174.900 93.700 175.000 ;
        RECT 94.200 174.800 94.600 175.000 ;
        RECT 95.800 174.800 96.200 175.000 ;
        RECT 104.600 174.700 105.000 175.000 ;
        RECT 92.600 174.100 97.000 174.500 ;
        RECT 97.300 174.300 98.300 174.700 ;
        RECT 100.200 174.300 101.800 174.700 ;
        RECT 77.300 172.700 77.700 172.800 ;
        RECT 74.200 172.100 74.600 172.500 ;
        RECT 76.300 172.400 77.700 172.700 ;
        RECT 78.200 172.400 78.600 172.800 ;
        RECT 76.300 172.100 76.600 172.400 ;
        RECT 79.000 172.100 79.400 172.500 ;
        RECT 73.900 171.800 74.600 172.100 ;
        RECT 73.900 171.100 74.500 171.800 ;
        RECT 76.200 171.100 76.600 172.100 ;
        RECT 78.400 171.800 79.400 172.100 ;
        RECT 78.400 171.100 78.800 171.800 ;
        RECT 80.600 171.100 81.000 173.500 ;
        RECT 82.200 173.400 84.200 173.800 ;
        RECT 85.400 173.400 86.600 173.800 ;
        RECT 87.100 173.400 88.200 173.800 ;
        RECT 88.700 173.400 89.800 173.800 ;
        RECT 90.500 173.400 91.400 173.800 ;
        RECT 82.200 171.100 82.600 173.400 ;
        RECT 83.800 171.100 84.200 173.400 ;
        RECT 86.200 171.100 86.600 173.400 ;
        RECT 87.800 171.100 88.200 173.400 ;
        RECT 89.400 171.100 89.800 173.400 ;
        RECT 91.000 171.100 91.400 173.400 ;
        RECT 92.600 171.100 93.000 174.100 ;
        RECT 93.800 173.400 95.300 173.800 ;
        RECT 94.900 173.100 95.300 173.400 ;
        RECT 97.900 173.100 98.300 174.300 ;
        RECT 99.000 173.400 99.400 174.200 ;
        RECT 101.600 173.900 102.000 174.000 ;
        RECT 99.800 173.600 102.000 173.900 ;
        RECT 99.800 173.500 100.200 173.600 ;
        RECT 103.000 173.200 103.400 174.600 ;
        RECT 105.900 174.300 107.800 174.700 ;
        RECT 105.900 173.700 106.300 174.300 ;
        RECT 108.100 174.000 108.400 175.000 ;
        RECT 99.800 173.100 100.200 173.200 ;
        RECT 94.900 172.700 96.200 173.100 ;
        RECT 97.900 172.800 100.200 173.100 ;
        RECT 100.600 172.800 101.400 173.200 ;
        RECT 102.900 172.800 103.400 173.200 ;
        RECT 105.400 173.400 106.300 173.700 ;
        RECT 107.800 173.700 108.400 174.000 ;
        RECT 105.400 173.100 105.800 173.400 ;
        RECT 95.800 171.100 96.200 172.700 ;
        RECT 104.600 172.700 105.800 173.100 ;
        RECT 96.600 171.100 97.000 172.500 ;
        RECT 97.400 171.100 97.800 172.500 ;
        RECT 98.200 171.100 98.600 172.500 ;
        RECT 99.800 171.100 100.200 172.500 ;
        RECT 101.400 171.100 101.800 172.500 ;
        RECT 102.200 171.100 102.600 172.500 ;
        RECT 103.000 171.100 103.400 172.500 ;
        RECT 103.800 171.100 104.200 172.500 ;
        RECT 104.600 171.100 105.000 172.700 ;
        RECT 107.800 171.100 108.200 173.700 ;
        RECT 108.700 173.400 109.100 175.600 ;
        RECT 111.800 174.800 112.300 175.200 ;
        RECT 111.900 174.400 112.300 174.800 ;
        RECT 112.800 174.900 113.100 175.900 ;
        RECT 112.800 174.500 113.300 174.900 ;
        RECT 112.800 173.700 113.100 174.500 ;
        RECT 113.600 174.200 113.900 175.900 ;
        RECT 115.800 175.600 116.200 179.900 ;
        RECT 117.400 175.600 117.800 179.900 ;
        RECT 119.000 175.600 119.400 179.900 ;
        RECT 120.600 175.600 121.000 179.900 ;
        RECT 123.500 176.300 123.900 179.900 ;
        RECT 123.000 175.900 123.900 176.300 ;
        RECT 115.000 175.200 116.200 175.600 ;
        RECT 116.700 175.200 117.800 175.600 ;
        RECT 118.300 175.200 119.400 175.600 ;
        RECT 120.100 175.200 121.000 175.600 ;
        RECT 113.400 174.100 113.900 174.200 ;
        RECT 114.200 174.800 114.600 175.200 ;
        RECT 114.200 174.100 114.500 174.800 ;
        RECT 113.400 173.800 114.500 174.100 ;
        RECT 115.000 173.800 115.400 175.200 ;
        RECT 116.700 174.500 117.100 175.200 ;
        RECT 118.300 174.500 118.700 175.200 ;
        RECT 120.100 174.500 120.500 175.200 ;
        RECT 115.800 174.100 117.100 174.500 ;
        RECT 117.500 174.100 118.700 174.500 ;
        RECT 119.200 174.100 120.500 174.500 ;
        RECT 123.100 174.200 123.400 175.900 ;
        RECT 123.800 175.100 124.200 175.600 ;
        RECT 124.600 175.100 125.000 179.900 ;
        RECT 126.500 176.300 126.900 179.900 ;
        RECT 126.500 175.900 127.400 176.300 ;
        RECT 126.200 175.100 126.600 175.600 ;
        RECT 123.800 174.800 126.600 175.100 ;
        RECT 116.700 173.800 117.100 174.100 ;
        RECT 118.300 173.800 118.700 174.100 ;
        RECT 120.100 173.800 120.500 174.100 ;
        RECT 123.000 173.800 123.400 174.200 ;
        RECT 108.600 173.100 109.100 173.400 ;
        RECT 111.800 173.400 113.100 173.700 ;
        RECT 109.400 173.100 109.800 173.200 ;
        RECT 108.600 172.800 109.800 173.100 ;
        RECT 108.600 171.100 109.000 172.800 ;
        RECT 111.800 171.100 112.200 173.400 ;
        RECT 113.600 173.100 113.900 173.800 ;
        RECT 115.000 173.400 116.200 173.800 ;
        RECT 116.700 173.400 117.800 173.800 ;
        RECT 118.300 173.400 119.400 173.800 ;
        RECT 120.100 173.400 121.000 173.800 ;
        RECT 113.400 172.800 113.900 173.100 ;
        RECT 113.400 171.100 113.800 172.800 ;
        RECT 115.800 171.100 116.200 173.400 ;
        RECT 117.400 171.100 117.800 173.400 ;
        RECT 119.000 171.100 119.400 173.400 ;
        RECT 120.600 171.100 121.000 173.400 ;
        RECT 122.200 172.400 122.600 173.200 ;
        RECT 123.100 172.200 123.400 173.800 ;
        RECT 123.000 171.100 123.400 172.200 ;
        RECT 124.600 171.100 125.000 174.800 ;
        RECT 127.000 174.200 127.300 175.900 ;
        RECT 127.000 173.800 127.400 174.200 ;
        RECT 125.400 172.400 125.800 173.200 ;
        RECT 127.000 172.200 127.300 173.800 ;
        RECT 127.800 173.100 128.200 173.200 ;
        RECT 128.600 173.100 129.000 179.900 ;
        RECT 131.000 176.000 131.400 179.900 ;
        RECT 132.600 177.600 133.000 179.900 ;
        RECT 130.900 175.600 131.400 176.000 ;
        RECT 131.700 177.300 133.000 177.600 ;
        RECT 131.700 176.500 132.000 177.300 ;
        RECT 134.200 177.200 134.600 179.900 ;
        RECT 135.800 178.500 136.200 179.900 ;
        RECT 136.600 178.500 137.000 179.900 ;
        RECT 137.400 178.500 137.800 179.900 ;
        RECT 134.900 177.200 137.000 177.600 ;
        RECT 133.300 176.800 134.600 177.200 ;
        RECT 138.200 176.800 138.600 179.900 ;
        RECT 139.800 177.500 140.200 179.900 ;
        RECT 141.400 177.500 141.800 179.900 ;
        RECT 142.200 178.500 142.600 179.900 ;
        RECT 143.000 178.500 143.400 179.900 ;
        RECT 144.600 177.600 145.000 179.900 ;
        RECT 146.200 178.200 146.600 179.900 ;
        RECT 150.200 178.200 150.600 179.900 ;
        RECT 146.200 177.900 146.700 178.200 ;
        RECT 146.400 177.600 146.700 177.900 ;
        RECT 150.100 177.900 150.600 178.200 ;
        RECT 150.100 177.600 150.400 177.900 ;
        RECT 151.800 177.600 152.200 179.900 ;
        RECT 153.400 178.500 153.800 179.900 ;
        RECT 154.200 178.500 154.600 179.900 ;
        RECT 144.000 177.200 146.100 177.600 ;
        RECT 146.400 177.300 147.400 177.600 ;
        RECT 139.800 176.800 141.100 177.200 ;
        RECT 141.400 176.900 144.300 177.200 ;
        RECT 145.800 177.000 146.100 177.200 ;
        RECT 135.800 176.500 136.200 176.600 ;
        RECT 131.700 176.200 136.200 176.500 ;
        RECT 137.400 176.500 137.800 176.600 ;
        RECT 141.400 176.500 141.700 176.900 ;
        RECT 144.600 176.600 145.300 176.900 ;
        RECT 145.800 176.600 146.600 177.000 ;
        RECT 137.400 176.200 141.700 176.500 ;
        RECT 142.200 176.500 145.300 176.600 ;
        RECT 142.200 176.300 144.900 176.500 ;
        RECT 142.200 176.200 142.600 176.300 ;
        RECT 129.400 174.100 129.800 174.200 ;
        RECT 130.900 174.100 131.300 175.600 ;
        RECT 131.700 175.300 132.000 176.200 ;
        RECT 129.400 173.800 131.300 174.100 ;
        RECT 129.400 173.400 129.800 173.800 ;
        RECT 130.900 173.400 131.300 173.800 ;
        RECT 131.600 175.000 132.000 175.300 ;
        RECT 135.000 175.000 146.700 175.300 ;
        RECT 131.600 174.000 131.900 175.000 ;
        RECT 135.000 174.700 135.400 175.000 ;
        RECT 143.800 174.800 144.200 175.000 ;
        RECT 146.200 174.900 146.700 175.000 ;
        RECT 146.200 174.800 146.600 174.900 ;
        RECT 132.200 174.300 134.100 174.700 ;
        RECT 131.600 173.700 132.200 174.000 ;
        RECT 127.800 172.800 129.000 173.100 ;
        RECT 130.900 173.000 131.400 173.400 ;
        RECT 127.800 172.400 128.200 172.800 ;
        RECT 127.000 171.100 127.400 172.200 ;
        RECT 128.600 171.100 129.000 172.800 ;
        RECT 131.000 171.100 131.400 173.000 ;
        RECT 131.800 171.100 132.200 173.700 ;
        RECT 133.700 173.700 134.100 174.300 ;
        RECT 133.700 173.400 134.600 173.700 ;
        RECT 134.200 173.100 134.600 173.400 ;
        RECT 136.600 173.200 137.000 174.600 ;
        RECT 138.200 174.300 139.800 174.700 ;
        RECT 141.700 174.300 142.700 174.700 ;
        RECT 147.000 174.500 147.400 177.300 ;
        RECT 138.000 173.900 138.400 174.000 ;
        RECT 138.000 173.600 140.200 173.900 ;
        RECT 139.800 173.500 140.200 173.600 ;
        RECT 140.600 173.400 141.000 174.200 ;
        RECT 134.200 172.700 135.400 173.100 ;
        RECT 136.600 172.800 137.100 173.200 ;
        RECT 138.600 172.800 139.400 173.200 ;
        RECT 139.800 173.100 140.200 173.200 ;
        RECT 141.700 173.100 142.100 174.300 ;
        RECT 143.000 174.100 147.400 174.500 ;
        RECT 144.700 173.400 146.200 173.800 ;
        RECT 144.700 173.100 145.100 173.400 ;
        RECT 139.800 172.800 142.100 173.100 ;
        RECT 135.000 171.100 135.400 172.700 ;
        RECT 143.800 172.700 145.100 173.100 ;
        RECT 135.800 171.100 136.200 172.500 ;
        RECT 136.600 171.100 137.000 172.500 ;
        RECT 137.400 171.100 137.800 172.500 ;
        RECT 138.200 171.100 138.600 172.500 ;
        RECT 139.800 171.100 140.200 172.500 ;
        RECT 141.400 171.100 141.800 172.500 ;
        RECT 142.200 171.100 142.600 172.500 ;
        RECT 143.000 171.100 143.400 172.500 ;
        RECT 143.800 171.100 144.200 172.700 ;
        RECT 147.000 171.100 147.400 174.100 ;
        RECT 149.400 177.300 150.400 177.600 ;
        RECT 149.400 174.500 149.800 177.300 ;
        RECT 150.700 177.200 152.800 177.600 ;
        RECT 155.000 177.500 155.400 179.900 ;
        RECT 156.600 177.500 157.000 179.900 ;
        RECT 150.700 177.000 151.000 177.200 ;
        RECT 150.200 176.600 151.000 177.000 ;
        RECT 152.500 176.900 155.400 177.200 ;
        RECT 151.500 176.600 152.200 176.900 ;
        RECT 151.500 176.500 154.600 176.600 ;
        RECT 151.900 176.300 154.600 176.500 ;
        RECT 154.200 176.200 154.600 176.300 ;
        RECT 155.100 176.500 155.400 176.900 ;
        RECT 155.700 176.800 157.000 177.200 ;
        RECT 158.200 176.800 158.600 179.900 ;
        RECT 159.000 178.500 159.400 179.900 ;
        RECT 159.800 178.500 160.200 179.900 ;
        RECT 160.600 178.500 161.000 179.900 ;
        RECT 159.800 177.200 161.900 177.600 ;
        RECT 162.200 177.200 162.600 179.900 ;
        RECT 163.800 177.600 164.200 179.900 ;
        RECT 163.800 177.300 165.100 177.600 ;
        RECT 162.200 176.800 163.500 177.200 ;
        RECT 159.000 176.500 159.400 176.600 ;
        RECT 155.100 176.200 159.400 176.500 ;
        RECT 160.600 176.500 161.000 176.600 ;
        RECT 164.800 176.500 165.100 177.300 ;
        RECT 160.600 176.200 165.100 176.500 ;
        RECT 164.800 175.300 165.100 176.200 ;
        RECT 165.400 176.000 165.800 179.900 ;
        RECT 165.400 175.600 165.900 176.000 ;
        RECT 150.100 175.000 161.800 175.300 ;
        RECT 164.800 175.000 165.200 175.300 ;
        RECT 150.100 174.900 150.500 175.000 ;
        RECT 151.000 174.800 151.400 175.000 ;
        RECT 152.600 174.800 153.000 175.000 ;
        RECT 161.400 174.700 161.800 175.000 ;
        RECT 149.400 174.100 153.800 174.500 ;
        RECT 154.100 174.300 155.100 174.700 ;
        RECT 157.000 174.300 158.600 174.700 ;
        RECT 149.400 171.100 149.800 174.100 ;
        RECT 150.600 173.400 152.100 173.800 ;
        RECT 151.700 173.100 152.100 173.400 ;
        RECT 154.700 173.100 155.100 174.300 ;
        RECT 155.800 173.400 156.200 174.200 ;
        RECT 158.400 173.900 158.800 174.000 ;
        RECT 156.600 173.600 158.800 173.900 ;
        RECT 156.600 173.500 157.000 173.600 ;
        RECT 159.800 173.200 160.200 174.600 ;
        RECT 162.700 174.300 164.600 174.700 ;
        RECT 162.700 173.700 163.100 174.300 ;
        RECT 164.900 174.000 165.200 175.000 ;
        RECT 156.600 173.100 157.000 173.200 ;
        RECT 151.700 172.700 153.000 173.100 ;
        RECT 154.700 172.800 157.000 173.100 ;
        RECT 157.400 172.800 158.200 173.200 ;
        RECT 159.700 172.800 160.200 173.200 ;
        RECT 162.200 173.400 163.100 173.700 ;
        RECT 164.600 173.700 165.200 174.000 ;
        RECT 162.200 173.100 162.600 173.400 ;
        RECT 152.600 171.100 153.000 172.700 ;
        RECT 161.400 172.700 162.600 173.100 ;
        RECT 153.400 171.100 153.800 172.500 ;
        RECT 154.200 171.100 154.600 172.500 ;
        RECT 155.000 171.100 155.400 172.500 ;
        RECT 156.600 171.100 157.000 172.500 ;
        RECT 158.200 171.100 158.600 172.500 ;
        RECT 159.000 171.100 159.400 172.500 ;
        RECT 159.800 171.100 160.200 172.500 ;
        RECT 160.600 171.100 161.000 172.500 ;
        RECT 161.400 171.100 161.800 172.700 ;
        RECT 164.600 171.100 165.000 173.700 ;
        RECT 165.500 173.400 165.900 175.600 ;
        RECT 167.800 175.600 168.200 179.900 ;
        RECT 169.400 175.600 169.800 179.900 ;
        RECT 171.000 175.600 171.400 179.900 ;
        RECT 172.600 175.600 173.000 179.900 ;
        RECT 175.000 178.200 175.400 179.900 ;
        RECT 174.900 177.900 175.400 178.200 ;
        RECT 174.900 177.600 175.200 177.900 ;
        RECT 176.600 177.600 177.000 179.900 ;
        RECT 178.200 178.500 178.600 179.900 ;
        RECT 179.000 178.500 179.400 179.900 ;
        RECT 174.200 177.300 175.200 177.600 ;
        RECT 167.800 175.200 168.700 175.600 ;
        RECT 169.400 175.200 170.500 175.600 ;
        RECT 171.000 175.200 172.100 175.600 ;
        RECT 172.600 175.200 173.800 175.600 ;
        RECT 168.300 174.500 168.700 175.200 ;
        RECT 170.100 174.500 170.500 175.200 ;
        RECT 171.700 174.500 172.100 175.200 ;
        RECT 168.300 174.100 169.600 174.500 ;
        RECT 170.100 174.100 171.300 174.500 ;
        RECT 171.700 174.100 173.000 174.500 ;
        RECT 168.300 173.800 168.700 174.100 ;
        RECT 170.100 173.800 170.500 174.100 ;
        RECT 171.700 173.800 172.100 174.100 ;
        RECT 173.400 173.800 173.800 175.200 ;
        RECT 165.400 173.000 165.900 173.400 ;
        RECT 167.800 173.400 168.700 173.800 ;
        RECT 169.400 173.400 170.500 173.800 ;
        RECT 171.000 173.400 172.100 173.800 ;
        RECT 172.600 173.400 173.800 173.800 ;
        RECT 174.200 174.500 174.600 177.300 ;
        RECT 175.500 177.200 177.600 177.600 ;
        RECT 179.800 177.500 180.200 179.900 ;
        RECT 181.400 177.500 181.800 179.900 ;
        RECT 175.500 177.000 175.800 177.200 ;
        RECT 175.000 176.600 175.800 177.000 ;
        RECT 177.300 176.900 180.200 177.200 ;
        RECT 176.300 176.600 177.000 176.900 ;
        RECT 176.300 176.500 179.400 176.600 ;
        RECT 176.700 176.300 179.400 176.500 ;
        RECT 179.000 176.200 179.400 176.300 ;
        RECT 179.900 176.500 180.200 176.900 ;
        RECT 180.500 176.800 181.800 177.200 ;
        RECT 183.000 176.800 183.400 179.900 ;
        RECT 183.800 178.500 184.200 179.900 ;
        RECT 184.600 178.500 185.000 179.900 ;
        RECT 185.400 178.500 185.800 179.900 ;
        RECT 184.600 177.200 186.700 177.600 ;
        RECT 187.000 177.200 187.400 179.900 ;
        RECT 188.600 177.600 189.000 179.900 ;
        RECT 188.600 177.300 189.900 177.600 ;
        RECT 187.000 176.800 188.300 177.200 ;
        RECT 183.800 176.500 184.200 176.600 ;
        RECT 179.900 176.200 184.200 176.500 ;
        RECT 185.400 176.500 185.800 176.600 ;
        RECT 189.600 176.500 189.900 177.300 ;
        RECT 185.400 176.200 189.900 176.500 ;
        RECT 189.600 175.300 189.900 176.200 ;
        RECT 190.200 176.000 190.600 179.900 ;
        RECT 190.200 175.600 190.700 176.000 ;
        RECT 174.900 175.000 186.600 175.300 ;
        RECT 189.600 175.000 190.000 175.300 ;
        RECT 174.900 174.900 175.300 175.000 ;
        RECT 177.400 174.800 177.800 175.000 ;
        RECT 186.200 174.700 186.600 175.000 ;
        RECT 174.200 174.100 178.600 174.500 ;
        RECT 178.900 174.300 179.900 174.700 ;
        RECT 181.800 174.300 183.400 174.700 ;
        RECT 165.400 171.100 165.800 173.000 ;
        RECT 167.800 171.100 168.200 173.400 ;
        RECT 169.400 171.100 169.800 173.400 ;
        RECT 171.000 171.100 171.400 173.400 ;
        RECT 172.600 171.100 173.000 173.400 ;
        RECT 174.200 171.100 174.600 174.100 ;
        RECT 175.400 173.400 176.900 173.800 ;
        RECT 176.500 173.100 176.900 173.400 ;
        RECT 179.500 173.100 179.900 174.300 ;
        RECT 180.600 173.400 181.000 174.200 ;
        RECT 183.200 173.900 183.600 174.000 ;
        RECT 181.400 173.600 183.600 173.900 ;
        RECT 181.400 173.500 181.800 173.600 ;
        RECT 184.600 173.200 185.000 174.600 ;
        RECT 187.500 174.300 189.400 174.700 ;
        RECT 187.500 173.700 187.900 174.300 ;
        RECT 189.700 174.000 190.000 175.000 ;
        RECT 181.400 173.100 181.800 173.200 ;
        RECT 176.500 172.700 177.800 173.100 ;
        RECT 179.500 172.800 181.800 173.100 ;
        RECT 182.200 172.800 183.000 173.200 ;
        RECT 184.500 172.800 185.000 173.200 ;
        RECT 187.000 173.400 187.900 173.700 ;
        RECT 189.400 173.700 190.000 174.000 ;
        RECT 187.000 173.100 187.400 173.400 ;
        RECT 177.400 171.100 177.800 172.700 ;
        RECT 186.200 172.700 187.400 173.100 ;
        RECT 178.200 171.100 178.600 172.500 ;
        RECT 179.000 171.100 179.400 172.500 ;
        RECT 179.800 171.100 180.200 172.500 ;
        RECT 181.400 171.100 181.800 172.500 ;
        RECT 183.000 171.100 183.400 172.500 ;
        RECT 183.800 171.100 184.200 172.500 ;
        RECT 184.600 171.100 185.000 172.500 ;
        RECT 185.400 171.100 185.800 172.500 ;
        RECT 186.200 171.100 186.600 172.700 ;
        RECT 189.400 171.100 189.800 173.700 ;
        RECT 190.300 173.400 190.700 175.600 ;
        RECT 190.200 173.000 190.700 173.400 ;
        RECT 190.200 171.100 190.600 173.000 ;
        RECT 191.800 171.100 192.200 179.900 ;
        RECT 194.200 177.900 194.600 179.900 ;
        RECT 194.300 177.800 194.600 177.900 ;
        RECT 195.800 177.900 196.200 179.900 ;
        RECT 195.800 177.800 196.100 177.900 ;
        RECT 194.300 177.500 196.100 177.800 ;
        RECT 195.000 176.400 195.400 177.200 ;
        RECT 195.800 176.200 196.100 177.500 ;
        RECT 195.800 175.800 196.200 176.200 ;
        RECT 194.200 174.800 195.000 175.200 ;
        RECT 195.800 174.200 196.100 175.800 ;
        RECT 195.300 174.100 196.100 174.200 ;
        RECT 195.200 173.900 196.100 174.100 ;
        RECT 197.400 175.100 197.800 179.900 ;
        RECT 198.200 176.200 198.600 179.900 ;
        RECT 198.200 175.900 199.300 176.200 ;
        RECT 199.000 175.600 199.300 175.900 ;
        RECT 199.000 175.200 199.600 175.600 ;
        RECT 198.200 175.100 198.600 175.200 ;
        RECT 197.400 174.800 198.600 175.100 ;
        RECT 195.200 173.200 195.600 173.900 ;
        RECT 192.600 172.400 193.000 173.200 ;
        RECT 195.000 172.800 195.600 173.200 ;
        RECT 195.200 171.100 195.600 172.800 ;
        RECT 196.600 172.400 197.000 173.200 ;
        RECT 197.400 171.100 197.800 174.800 ;
        RECT 198.200 174.400 198.600 174.800 ;
        RECT 199.000 173.700 199.300 175.200 ;
        RECT 198.200 173.400 199.300 173.700 ;
        RECT 201.400 175.100 201.800 179.900 ;
        RECT 202.200 176.200 202.600 179.900 ;
        RECT 202.200 175.900 203.300 176.200 ;
        RECT 203.000 175.600 203.300 175.900 ;
        RECT 203.000 175.200 203.600 175.600 ;
        RECT 202.200 175.100 202.600 175.200 ;
        RECT 201.400 174.800 202.600 175.100 ;
        RECT 198.200 171.100 198.600 173.400 ;
        RECT 200.600 172.400 201.000 173.200 ;
        RECT 201.400 171.100 201.800 174.800 ;
        RECT 202.200 174.400 202.600 174.800 ;
        RECT 203.000 173.700 203.300 175.200 ;
        RECT 202.200 173.400 203.300 173.700 ;
        RECT 202.200 171.100 202.600 173.400 ;
        RECT 1.400 168.000 1.800 169.900 ;
        RECT 1.300 167.600 1.800 168.000 ;
        RECT 1.300 165.400 1.700 167.600 ;
        RECT 2.200 167.300 2.600 169.900 ;
        RECT 5.400 168.300 5.800 169.900 ;
        RECT 6.200 168.500 6.600 169.900 ;
        RECT 7.000 168.500 7.400 169.900 ;
        RECT 7.800 168.500 8.200 169.900 ;
        RECT 8.600 168.500 9.000 169.900 ;
        RECT 10.200 168.500 10.600 169.900 ;
        RECT 11.800 168.500 12.200 169.900 ;
        RECT 12.600 168.500 13.000 169.900 ;
        RECT 13.400 168.500 13.800 169.900 ;
        RECT 4.600 167.900 5.800 168.300 ;
        RECT 14.200 168.300 14.600 169.900 ;
        RECT 4.600 167.600 5.000 167.900 ;
        RECT 2.000 167.000 2.600 167.300 ;
        RECT 4.100 167.300 5.000 167.600 ;
        RECT 7.000 167.800 7.500 168.200 ;
        RECT 9.000 167.800 9.800 168.200 ;
        RECT 10.200 167.900 12.500 168.200 ;
        RECT 14.200 167.900 15.500 168.300 ;
        RECT 10.200 167.800 10.600 167.900 ;
        RECT 2.000 166.000 2.300 167.000 ;
        RECT 4.100 166.700 4.500 167.300 ;
        RECT 2.600 166.300 4.500 166.700 ;
        RECT 7.000 166.400 7.400 167.800 ;
        RECT 10.200 167.400 10.600 167.500 ;
        RECT 8.400 167.100 10.600 167.400 ;
        RECT 8.400 167.000 8.800 167.100 ;
        RECT 11.000 166.800 11.400 167.600 ;
        RECT 12.100 166.700 12.500 167.900 ;
        RECT 15.100 167.600 15.500 167.900 ;
        RECT 15.100 167.200 16.600 167.600 ;
        RECT 17.400 166.900 17.800 169.900 ;
        RECT 19.000 168.000 19.400 169.900 ;
        RECT 8.600 166.300 10.200 166.700 ;
        RECT 12.100 166.300 13.100 166.700 ;
        RECT 13.400 166.500 17.800 166.900 ;
        RECT 5.400 166.000 5.800 166.300 ;
        RECT 14.200 166.000 14.600 166.200 ;
        RECT 15.800 166.000 16.200 166.200 ;
        RECT 16.700 166.000 17.100 166.100 ;
        RECT 2.000 165.700 2.400 166.000 ;
        RECT 5.400 165.700 17.100 166.000 ;
        RECT 1.300 165.000 1.800 165.400 ;
        RECT 1.400 161.100 1.800 165.000 ;
        RECT 2.100 164.800 2.400 165.700 ;
        RECT 2.100 164.500 6.600 164.800 ;
        RECT 2.100 163.700 2.400 164.500 ;
        RECT 6.200 164.400 6.600 164.500 ;
        RECT 7.800 164.500 12.100 164.800 ;
        RECT 7.800 164.400 8.200 164.500 ;
        RECT 3.700 163.800 5.000 164.200 ;
        RECT 2.100 163.400 3.400 163.700 ;
        RECT 3.000 161.100 3.400 163.400 ;
        RECT 4.600 161.100 5.000 163.800 ;
        RECT 5.300 163.400 7.400 163.800 ;
        RECT 6.200 161.100 6.600 162.500 ;
        RECT 7.000 161.100 7.400 162.500 ;
        RECT 7.800 161.100 8.200 162.500 ;
        RECT 8.600 161.100 9.000 164.200 ;
        RECT 10.200 163.800 11.500 164.200 ;
        RECT 11.800 164.100 12.100 164.500 ;
        RECT 12.600 164.700 13.000 164.800 ;
        RECT 12.600 164.500 15.300 164.700 ;
        RECT 12.600 164.400 15.700 164.500 ;
        RECT 15.000 164.100 15.700 164.400 ;
        RECT 11.800 163.800 14.700 164.100 ;
        RECT 16.200 164.000 17.000 164.400 ;
        RECT 16.200 163.800 16.500 164.000 ;
        RECT 10.200 161.100 10.600 163.500 ;
        RECT 11.800 161.100 12.200 163.500 ;
        RECT 14.400 163.400 16.500 163.800 ;
        RECT 17.400 163.700 17.800 166.500 ;
        RECT 18.900 167.600 19.400 168.000 ;
        RECT 18.900 165.400 19.300 167.600 ;
        RECT 19.800 167.300 20.200 169.900 ;
        RECT 23.000 168.300 23.400 169.900 ;
        RECT 23.800 168.500 24.200 169.900 ;
        RECT 24.600 168.500 25.000 169.900 ;
        RECT 25.400 168.500 25.800 169.900 ;
        RECT 26.200 168.500 26.600 169.900 ;
        RECT 27.800 168.500 28.200 169.900 ;
        RECT 29.400 168.500 29.800 169.900 ;
        RECT 30.200 168.500 30.600 169.900 ;
        RECT 31.000 168.500 31.400 169.900 ;
        RECT 22.200 167.900 23.400 168.300 ;
        RECT 31.800 168.300 32.200 169.900 ;
        RECT 22.200 167.600 22.600 167.900 ;
        RECT 19.600 167.000 20.200 167.300 ;
        RECT 21.700 167.300 22.600 167.600 ;
        RECT 24.600 167.800 25.100 168.200 ;
        RECT 26.600 167.800 27.400 168.200 ;
        RECT 27.800 167.900 30.100 168.200 ;
        RECT 31.800 167.900 33.100 168.300 ;
        RECT 27.800 167.800 28.200 167.900 ;
        RECT 19.600 166.000 19.900 167.000 ;
        RECT 21.700 166.700 22.100 167.300 ;
        RECT 20.200 166.300 22.100 166.700 ;
        RECT 23.000 166.800 23.400 167.200 ;
        RECT 23.000 166.300 23.300 166.800 ;
        RECT 24.600 166.400 25.000 167.800 ;
        RECT 27.800 167.400 28.200 167.500 ;
        RECT 26.000 167.100 28.200 167.400 ;
        RECT 26.000 167.000 26.400 167.100 ;
        RECT 28.600 166.800 29.000 167.600 ;
        RECT 29.700 166.700 30.100 167.900 ;
        RECT 32.700 167.600 33.100 167.900 ;
        RECT 32.700 167.200 34.200 167.600 ;
        RECT 35.000 166.900 35.400 169.900 ;
        RECT 36.600 168.000 37.000 169.900 ;
        RECT 26.200 166.300 27.800 166.700 ;
        RECT 29.700 166.300 30.700 166.700 ;
        RECT 31.000 166.500 35.400 166.900 ;
        RECT 23.000 166.000 23.400 166.300 ;
        RECT 31.800 166.000 32.200 166.200 ;
        RECT 33.400 166.000 33.800 166.200 ;
        RECT 34.300 166.000 34.700 166.100 ;
        RECT 19.600 165.700 20.000 166.000 ;
        RECT 23.000 165.700 34.700 166.000 ;
        RECT 18.900 165.000 19.400 165.400 ;
        RECT 16.800 163.400 17.800 163.700 ;
        RECT 12.600 161.100 13.000 162.500 ;
        RECT 13.400 161.100 13.800 162.500 ;
        RECT 15.000 161.100 15.400 163.400 ;
        RECT 16.800 163.100 17.100 163.400 ;
        RECT 16.600 162.800 17.100 163.100 ;
        RECT 16.600 161.100 17.000 162.800 ;
        RECT 19.000 161.100 19.400 165.000 ;
        RECT 19.700 164.800 20.000 165.700 ;
        RECT 19.700 164.500 24.200 164.800 ;
        RECT 19.700 163.700 20.000 164.500 ;
        RECT 23.800 164.400 24.200 164.500 ;
        RECT 25.400 164.500 29.700 164.800 ;
        RECT 25.400 164.400 25.800 164.500 ;
        RECT 21.300 163.800 22.600 164.200 ;
        RECT 19.700 163.400 21.000 163.700 ;
        RECT 20.600 161.100 21.000 163.400 ;
        RECT 22.200 161.100 22.600 163.800 ;
        RECT 22.900 163.400 25.000 163.800 ;
        RECT 23.800 161.100 24.200 162.500 ;
        RECT 24.600 161.100 25.000 162.500 ;
        RECT 25.400 161.100 25.800 162.500 ;
        RECT 26.200 161.100 26.600 164.200 ;
        RECT 27.800 163.800 29.100 164.200 ;
        RECT 29.400 164.100 29.700 164.500 ;
        RECT 30.200 164.700 30.600 164.800 ;
        RECT 30.200 164.500 32.900 164.700 ;
        RECT 30.200 164.400 33.300 164.500 ;
        RECT 32.600 164.100 33.300 164.400 ;
        RECT 29.400 163.800 32.300 164.100 ;
        RECT 33.800 164.000 34.600 164.400 ;
        RECT 33.800 163.800 34.100 164.000 ;
        RECT 27.800 161.100 28.200 163.500 ;
        RECT 29.400 161.100 29.800 163.500 ;
        RECT 32.000 163.400 34.100 163.800 ;
        RECT 35.000 163.700 35.400 166.500 ;
        RECT 36.500 167.600 37.000 168.000 ;
        RECT 36.500 165.400 36.900 167.600 ;
        RECT 37.400 167.300 37.800 169.900 ;
        RECT 40.600 168.300 41.000 169.900 ;
        RECT 41.400 168.500 41.800 169.900 ;
        RECT 42.200 168.500 42.600 169.900 ;
        RECT 43.000 168.500 43.400 169.900 ;
        RECT 43.800 168.500 44.200 169.900 ;
        RECT 45.400 168.500 45.800 169.900 ;
        RECT 47.000 168.500 47.400 169.900 ;
        RECT 47.800 168.500 48.200 169.900 ;
        RECT 48.600 168.500 49.000 169.900 ;
        RECT 39.800 167.900 41.000 168.300 ;
        RECT 49.400 168.300 49.800 169.900 ;
        RECT 39.800 167.600 40.200 167.900 ;
        RECT 37.200 167.000 37.800 167.300 ;
        RECT 39.300 167.300 40.200 167.600 ;
        RECT 42.200 167.800 42.700 168.200 ;
        RECT 44.200 167.800 45.000 168.200 ;
        RECT 45.400 167.900 47.700 168.200 ;
        RECT 49.400 167.900 50.700 168.300 ;
        RECT 45.400 167.800 45.800 167.900 ;
        RECT 37.200 166.000 37.500 167.000 ;
        RECT 39.300 166.700 39.700 167.300 ;
        RECT 37.800 166.300 39.700 166.700 ;
        RECT 42.200 166.400 42.600 167.800 ;
        RECT 45.400 167.400 45.800 167.500 ;
        RECT 43.600 167.100 45.800 167.400 ;
        RECT 43.600 167.000 44.000 167.100 ;
        RECT 46.200 166.800 46.600 167.600 ;
        RECT 47.300 166.700 47.700 167.900 ;
        RECT 50.300 167.600 50.700 167.900 ;
        RECT 50.300 167.200 51.800 167.600 ;
        RECT 52.600 166.900 53.000 169.900 ;
        RECT 55.800 168.200 56.200 169.900 ;
        RECT 55.700 167.900 56.200 168.200 ;
        RECT 55.700 167.200 56.000 167.900 ;
        RECT 57.400 167.600 57.800 169.900 ;
        RECT 58.200 168.000 58.600 169.900 ;
        RECT 59.800 168.000 60.200 169.900 ;
        RECT 58.200 167.900 60.200 168.000 ;
        RECT 60.600 167.900 61.000 169.900 ;
        RECT 61.700 168.200 62.100 169.900 ;
        RECT 61.700 167.900 62.600 168.200 ;
        RECT 58.300 167.700 60.100 167.900 ;
        RECT 56.500 167.300 57.800 167.600 ;
        RECT 43.800 166.300 45.400 166.700 ;
        RECT 47.300 166.300 48.300 166.700 ;
        RECT 48.600 166.500 53.000 166.900 ;
        RECT 53.400 167.100 53.800 167.200 ;
        RECT 55.700 167.100 56.200 167.200 ;
        RECT 53.400 166.800 56.200 167.100 ;
        RECT 40.600 166.000 41.000 166.300 ;
        RECT 49.400 166.000 49.800 166.200 ;
        RECT 51.000 166.000 51.400 166.200 ;
        RECT 51.900 166.000 52.300 166.100 ;
        RECT 37.200 165.700 37.600 166.000 ;
        RECT 40.600 165.700 52.300 166.000 ;
        RECT 36.500 165.000 37.000 165.400 ;
        RECT 34.400 163.400 35.400 163.700 ;
        RECT 30.200 161.100 30.600 162.500 ;
        RECT 31.000 161.100 31.400 162.500 ;
        RECT 32.600 161.100 33.000 163.400 ;
        RECT 34.400 163.100 34.700 163.400 ;
        RECT 34.200 162.800 34.700 163.100 ;
        RECT 34.200 161.100 34.600 162.800 ;
        RECT 36.600 161.100 37.000 165.000 ;
        RECT 37.300 164.800 37.600 165.700 ;
        RECT 37.300 164.500 41.800 164.800 ;
        RECT 37.300 163.700 37.600 164.500 ;
        RECT 41.400 164.400 41.800 164.500 ;
        RECT 43.000 164.500 47.300 164.800 ;
        RECT 43.000 164.400 43.400 164.500 ;
        RECT 38.900 163.800 40.200 164.200 ;
        RECT 37.300 163.400 38.600 163.700 ;
        RECT 38.200 161.100 38.600 163.400 ;
        RECT 39.800 161.100 40.200 163.800 ;
        RECT 40.500 163.400 42.600 163.800 ;
        RECT 41.400 161.100 41.800 162.500 ;
        RECT 42.200 161.100 42.600 162.500 ;
        RECT 43.000 161.100 43.400 162.500 ;
        RECT 43.800 161.100 44.200 164.200 ;
        RECT 45.400 163.800 46.700 164.200 ;
        RECT 47.000 164.100 47.300 164.500 ;
        RECT 47.800 164.700 48.200 164.800 ;
        RECT 47.800 164.500 50.500 164.700 ;
        RECT 47.800 164.400 50.900 164.500 ;
        RECT 50.200 164.100 50.900 164.400 ;
        RECT 47.000 163.800 49.900 164.100 ;
        RECT 51.400 164.000 52.200 164.400 ;
        RECT 51.400 163.800 51.700 164.000 ;
        RECT 45.400 161.100 45.800 163.500 ;
        RECT 47.000 161.100 47.400 163.500 ;
        RECT 49.600 163.400 51.700 163.800 ;
        RECT 52.600 163.700 53.000 166.500 ;
        RECT 55.700 165.100 56.000 166.800 ;
        RECT 56.500 166.500 56.800 167.300 ;
        RECT 58.600 167.200 59.000 167.400 ;
        RECT 60.600 167.200 60.900 167.900 ;
        RECT 58.200 166.900 59.000 167.200 ;
        RECT 58.200 166.800 58.600 166.900 ;
        RECT 59.700 166.800 61.000 167.200 ;
        RECT 56.300 166.100 56.800 166.500 ;
        RECT 56.500 165.100 56.800 166.100 ;
        RECT 57.300 166.200 57.700 166.600 ;
        RECT 57.300 165.800 57.800 166.200 ;
        RECT 59.000 165.800 59.400 166.600 ;
        RECT 59.700 165.100 60.000 166.800 ;
        RECT 62.200 166.100 62.600 167.900 ;
        RECT 65.400 167.900 65.800 169.900 ;
        RECT 67.800 168.900 68.200 169.900 ;
        RECT 66.100 168.200 66.500 168.600 ;
        RECT 66.200 168.100 66.600 168.200 ;
        RECT 67.800 168.100 68.100 168.900 ;
        RECT 63.000 166.800 63.400 167.600 ;
        RECT 64.600 166.400 65.000 167.200 ;
        RECT 60.600 165.800 62.600 166.100 ;
        RECT 63.800 166.100 64.200 166.200 ;
        RECT 65.400 166.100 65.700 167.900 ;
        RECT 66.200 167.800 68.100 168.100 ;
        RECT 68.600 167.800 69.000 168.600 ;
        RECT 67.800 167.200 68.100 167.800 ;
        RECT 69.400 167.500 69.800 169.900 ;
        RECT 71.600 169.200 72.000 169.900 ;
        RECT 71.000 168.900 72.000 169.200 ;
        RECT 73.800 168.900 74.200 169.900 ;
        RECT 75.900 169.200 76.500 169.900 ;
        RECT 75.800 168.900 76.500 169.200 ;
        RECT 71.000 168.500 71.400 168.900 ;
        RECT 73.800 168.600 74.100 168.900 ;
        RECT 71.800 168.200 72.200 168.600 ;
        RECT 72.700 168.300 74.100 168.600 ;
        RECT 75.800 168.500 76.200 168.900 ;
        RECT 72.700 168.200 73.100 168.300 ;
        RECT 67.800 166.800 68.200 167.200 ;
        RECT 69.800 167.100 70.600 167.200 ;
        RECT 71.900 167.100 72.200 168.200 ;
        RECT 76.700 167.700 77.100 167.800 ;
        RECT 78.200 167.700 78.600 169.900 ;
        RECT 79.000 168.000 79.400 169.900 ;
        RECT 80.600 168.000 81.000 169.900 ;
        RECT 79.000 167.900 81.000 168.000 ;
        RECT 81.400 167.900 81.800 169.900 ;
        RECT 82.500 168.200 82.900 169.900 ;
        RECT 82.500 167.900 83.400 168.200 ;
        RECT 79.100 167.700 80.900 167.900 ;
        RECT 76.700 167.400 78.600 167.700 ;
        RECT 74.700 167.100 75.100 167.200 ;
        RECT 69.800 166.800 75.300 167.100 ;
        RECT 66.200 166.100 66.600 166.200 ;
        RECT 63.800 165.800 64.600 166.100 ;
        RECT 65.400 165.800 66.600 166.100 ;
        RECT 60.600 165.200 60.900 165.800 ;
        RECT 60.600 165.100 61.000 165.200 ;
        RECT 55.700 164.600 56.200 165.100 ;
        RECT 56.500 164.800 57.800 165.100 ;
        RECT 52.000 163.400 53.000 163.700 ;
        RECT 47.800 161.100 48.200 162.500 ;
        RECT 48.600 161.100 49.000 162.500 ;
        RECT 50.200 161.100 50.600 163.400 ;
        RECT 52.000 163.100 52.300 163.400 ;
        RECT 51.800 162.800 52.300 163.100 ;
        RECT 51.800 161.100 52.200 162.800 ;
        RECT 55.800 161.100 56.200 164.600 ;
        RECT 57.400 161.100 57.800 164.800 ;
        RECT 59.500 164.800 60.000 165.100 ;
        RECT 60.300 164.800 61.000 165.100 ;
        RECT 59.500 161.100 59.900 164.800 ;
        RECT 60.300 164.200 60.600 164.800 ;
        RECT 61.400 164.400 61.800 165.200 ;
        RECT 60.200 163.800 60.600 164.200 ;
        RECT 62.200 161.100 62.600 165.800 ;
        RECT 64.200 165.600 64.600 165.800 ;
        RECT 66.200 165.100 66.500 165.800 ;
        RECT 67.000 165.400 67.400 166.200 ;
        RECT 67.800 165.100 68.100 166.800 ;
        RECT 71.300 166.700 71.700 166.800 ;
        RECT 70.500 166.200 70.900 166.300 ;
        RECT 71.800 166.200 72.200 166.300 ;
        RECT 75.000 166.200 75.300 166.800 ;
        RECT 75.800 166.400 76.200 166.500 ;
        RECT 70.500 165.900 73.000 166.200 ;
        RECT 72.600 165.800 73.000 165.900 ;
        RECT 75.000 165.800 75.400 166.200 ;
        RECT 75.800 166.100 77.700 166.400 ;
        RECT 77.300 166.000 77.700 166.100 ;
        RECT 69.400 165.500 72.200 165.600 ;
        RECT 69.400 165.400 72.300 165.500 ;
        RECT 69.400 165.300 74.300 165.400 ;
        RECT 63.800 164.800 65.800 165.100 ;
        RECT 63.800 161.100 64.200 164.800 ;
        RECT 65.400 161.100 65.800 164.800 ;
        RECT 66.200 161.100 66.600 165.100 ;
        RECT 67.300 164.700 68.200 165.100 ;
        RECT 67.300 161.100 67.700 164.700 ;
        RECT 69.400 161.100 69.800 165.300 ;
        RECT 71.900 165.100 74.300 165.300 ;
        RECT 71.000 164.500 73.700 164.800 ;
        RECT 71.000 164.400 71.400 164.500 ;
        RECT 73.300 164.400 73.700 164.500 ;
        RECT 74.000 164.500 74.300 165.100 ;
        RECT 75.000 165.200 75.300 165.800 ;
        RECT 76.500 165.700 76.900 165.800 ;
        RECT 78.200 165.700 78.600 167.400 ;
        RECT 79.400 167.200 79.800 167.400 ;
        RECT 81.400 167.200 81.700 167.900 ;
        RECT 79.000 166.900 79.800 167.200 ;
        RECT 80.500 167.100 81.800 167.200 ;
        RECT 82.200 167.100 82.600 167.200 ;
        RECT 79.000 166.800 79.400 166.900 ;
        RECT 80.500 166.800 82.600 167.100 ;
        RECT 79.000 166.100 79.400 166.200 ;
        RECT 79.800 166.100 80.200 166.600 ;
        RECT 79.000 165.800 80.200 166.100 ;
        RECT 76.500 165.400 78.600 165.700 ;
        RECT 75.000 164.900 76.200 165.200 ;
        RECT 74.700 164.500 75.100 164.600 ;
        RECT 74.000 164.200 75.100 164.500 ;
        RECT 75.900 164.400 76.200 164.900 ;
        RECT 75.900 164.000 76.600 164.400 ;
        RECT 72.700 163.700 73.100 163.800 ;
        RECT 74.100 163.700 74.500 163.800 ;
        RECT 71.000 163.100 71.400 163.500 ;
        RECT 72.700 163.400 74.500 163.700 ;
        RECT 73.800 163.100 74.100 163.400 ;
        RECT 75.800 163.100 76.200 163.500 ;
        RECT 71.000 162.800 72.000 163.100 ;
        RECT 71.600 161.100 72.000 162.800 ;
        RECT 73.800 161.100 74.200 163.100 ;
        RECT 75.900 161.100 76.500 163.100 ;
        RECT 78.200 161.100 78.600 165.400 ;
        RECT 80.500 165.100 80.800 166.800 ;
        RECT 83.000 166.100 83.400 167.900 ;
        RECT 84.600 167.700 85.000 169.900 ;
        RECT 86.700 169.200 87.300 169.900 ;
        RECT 86.700 168.900 87.400 169.200 ;
        RECT 89.000 168.900 89.400 169.900 ;
        RECT 91.200 169.200 91.600 169.900 ;
        RECT 91.200 168.900 92.200 169.200 ;
        RECT 87.000 168.500 87.400 168.900 ;
        RECT 89.100 168.600 89.400 168.900 ;
        RECT 89.100 168.300 90.500 168.600 ;
        RECT 90.100 168.200 90.500 168.300 ;
        RECT 91.000 168.200 91.400 168.600 ;
        RECT 91.800 168.500 92.200 168.900 ;
        RECT 86.100 167.700 86.500 167.800 ;
        RECT 83.800 166.800 84.200 167.600 ;
        RECT 84.600 167.400 86.500 167.700 ;
        RECT 81.400 165.800 83.400 166.100 ;
        RECT 81.400 165.200 81.700 165.800 ;
        RECT 81.400 165.100 81.800 165.200 ;
        RECT 80.300 164.800 80.800 165.100 ;
        RECT 81.100 164.800 81.800 165.100 ;
        RECT 80.300 161.100 80.700 164.800 ;
        RECT 81.100 164.200 81.400 164.800 ;
        RECT 82.200 164.400 82.600 165.200 ;
        RECT 81.000 163.800 81.400 164.200 ;
        RECT 83.000 161.100 83.400 165.800 ;
        RECT 84.600 165.700 85.000 167.400 ;
        RECT 88.100 167.100 88.500 167.200 ;
        RECT 91.000 167.100 91.300 168.200 ;
        RECT 93.400 167.500 93.800 169.900 ;
        RECT 94.200 167.900 94.600 169.900 ;
        RECT 96.400 168.100 97.200 169.900 ;
        RECT 94.200 167.600 95.300 167.900 ;
        RECT 95.800 167.700 96.600 167.800 ;
        RECT 94.900 167.500 95.300 167.600 ;
        RECT 95.600 167.400 96.600 167.700 ;
        RECT 95.600 167.200 95.900 167.400 ;
        RECT 92.600 167.100 93.400 167.200 ;
        RECT 87.900 166.800 93.400 167.100 ;
        RECT 94.200 166.900 95.900 167.200 ;
        RECT 94.200 166.800 95.000 166.900 ;
        RECT 87.000 166.400 87.400 166.500 ;
        RECT 85.500 166.100 87.400 166.400 ;
        RECT 85.500 166.000 85.900 166.100 ;
        RECT 86.300 165.700 86.700 165.800 ;
        RECT 84.600 165.400 86.700 165.700 ;
        RECT 83.800 164.100 84.200 164.200 ;
        RECT 84.600 164.100 85.000 165.400 ;
        RECT 87.900 165.200 88.200 166.800 ;
        RECT 91.500 166.700 91.900 166.800 ;
        RECT 96.200 166.700 96.600 167.100 ;
        RECT 96.200 166.400 96.500 166.700 ;
        RECT 92.300 166.200 92.700 166.300 ;
        RECT 90.200 165.900 92.700 166.200 ;
        RECT 95.200 166.100 96.500 166.400 ;
        RECT 96.900 166.400 97.200 168.100 ;
        RECT 99.000 167.900 99.400 169.900 ;
        RECT 97.500 167.400 97.900 167.800 ;
        RECT 98.200 167.600 99.400 167.900 ;
        RECT 98.200 167.500 98.600 167.600 ;
        RECT 97.600 167.200 97.900 167.400 ;
        RECT 97.600 166.800 98.000 167.200 ;
        RECT 98.600 166.800 99.400 167.200 ;
        RECT 96.900 166.200 97.400 166.400 ;
        RECT 96.900 166.100 97.800 166.200 ;
        RECT 95.200 166.000 95.600 166.100 ;
        RECT 90.200 165.800 90.600 165.900 ;
        RECT 97.100 165.800 97.800 166.100 ;
        RECT 99.000 166.100 99.400 166.200 ;
        RECT 99.800 166.100 100.200 169.900 ;
        RECT 103.800 168.900 104.200 169.900 ;
        RECT 100.600 166.800 101.000 167.600 ;
        RECT 103.800 167.200 104.100 168.900 ;
        RECT 104.600 167.800 105.000 168.600 ;
        RECT 106.700 168.200 107.100 169.900 ;
        RECT 106.200 167.900 107.100 168.200 ;
        RECT 108.600 168.900 109.000 169.900 ;
        RECT 111.000 168.900 111.400 169.900 ;
        RECT 103.800 166.800 104.200 167.200 ;
        RECT 105.400 166.800 105.800 167.600 ;
        RECT 103.000 166.100 103.400 166.200 ;
        RECT 99.000 165.800 103.400 166.100 ;
        RECT 96.300 165.700 96.700 165.800 ;
        RECT 91.000 165.500 93.800 165.600 ;
        RECT 90.900 165.400 93.800 165.500 ;
        RECT 87.000 164.900 88.200 165.200 ;
        RECT 88.900 165.300 93.800 165.400 ;
        RECT 88.900 165.100 91.300 165.300 ;
        RECT 87.000 164.400 87.300 164.900 ;
        RECT 86.600 164.200 87.300 164.400 ;
        RECT 88.100 164.500 88.500 164.600 ;
        RECT 88.900 164.500 89.200 165.100 ;
        RECT 88.100 164.200 89.200 164.500 ;
        RECT 89.500 164.500 92.200 164.800 ;
        RECT 89.500 164.400 89.900 164.500 ;
        RECT 91.800 164.400 92.200 164.500 ;
        RECT 83.800 163.800 85.000 164.100 ;
        RECT 86.200 164.000 87.300 164.200 ;
        RECT 86.200 163.800 86.900 164.000 ;
        RECT 84.600 161.100 85.000 163.800 ;
        RECT 88.700 163.700 89.100 163.800 ;
        RECT 90.100 163.700 90.500 163.800 ;
        RECT 87.000 163.100 87.400 163.500 ;
        RECT 88.700 163.400 90.500 163.700 ;
        RECT 89.100 163.100 89.400 163.400 ;
        RECT 91.800 163.100 92.200 163.500 ;
        RECT 86.700 161.100 87.300 163.100 ;
        RECT 89.000 161.100 89.400 163.100 ;
        RECT 91.200 162.800 92.200 163.100 ;
        RECT 91.200 161.100 91.600 162.800 ;
        RECT 93.400 161.100 93.800 165.300 ;
        RECT 95.000 165.400 96.700 165.700 ;
        RECT 95.000 165.100 95.300 165.400 ;
        RECT 97.100 165.100 97.400 165.800 ;
        RECT 94.200 164.800 95.300 165.100 ;
        RECT 94.200 161.100 94.600 164.800 ;
        RECT 94.900 164.700 95.300 164.800 ;
        RECT 96.400 164.800 97.400 165.100 ;
        RECT 98.200 164.800 99.400 165.100 ;
        RECT 96.400 161.100 97.200 164.800 ;
        RECT 98.200 164.700 98.600 164.800 ;
        RECT 99.000 161.100 99.400 164.800 ;
        RECT 99.800 161.100 100.200 165.800 ;
        RECT 103.000 165.400 103.400 165.800 ;
        RECT 103.800 165.100 104.100 166.800 ;
        RECT 103.300 164.700 104.200 165.100 ;
        RECT 103.300 162.200 103.700 164.700 ;
        RECT 103.000 161.800 103.700 162.200 ;
        RECT 103.300 161.100 103.700 161.800 ;
        RECT 106.200 161.100 106.600 167.900 ;
        RECT 108.600 167.200 108.900 168.900 ;
        RECT 109.400 167.800 109.800 168.600 ;
        RECT 111.000 167.200 111.300 168.900 ;
        RECT 111.800 168.100 112.200 168.600 ;
        RECT 112.900 168.200 113.300 169.900 ;
        RECT 112.900 168.100 113.800 168.200 ;
        RECT 111.800 167.800 113.800 168.100 ;
        RECT 108.600 166.800 109.000 167.200 ;
        RECT 111.000 166.800 111.400 167.200 ;
        RECT 107.000 166.100 107.400 166.200 ;
        RECT 107.800 166.100 108.200 166.200 ;
        RECT 107.000 165.800 108.200 166.100 ;
        RECT 107.800 165.400 108.200 165.800 ;
        RECT 108.600 165.200 108.900 166.800 ;
        RECT 109.400 166.100 109.800 166.200 ;
        RECT 110.200 166.100 110.600 166.200 ;
        RECT 109.400 165.800 110.600 166.100 ;
        RECT 110.200 165.400 110.600 165.800 ;
        RECT 111.000 166.100 111.300 166.800 ;
        RECT 111.800 166.100 112.200 166.200 ;
        RECT 111.000 165.800 112.200 166.100 ;
        RECT 107.000 164.400 107.400 165.200 ;
        RECT 108.600 165.100 109.000 165.200 ;
        RECT 111.000 165.100 111.300 165.800 ;
        RECT 108.100 164.700 109.000 165.100 ;
        RECT 110.500 164.700 111.400 165.100 ;
        RECT 108.100 161.100 108.500 164.700 ;
        RECT 110.500 161.100 110.900 164.700 ;
        RECT 112.600 164.400 113.000 165.200 ;
        RECT 113.400 161.100 113.800 167.800 ;
        RECT 114.200 166.800 114.600 167.600 ;
        RECT 116.800 167.100 117.200 169.900 ;
        RECT 118.200 168.000 118.600 169.900 ;
        RECT 119.800 168.000 120.200 169.900 ;
        RECT 118.200 167.900 120.200 168.000 ;
        RECT 120.600 167.900 121.000 169.900 ;
        RECT 122.200 168.900 122.600 169.900 ;
        RECT 124.600 168.900 125.000 169.900 ;
        RECT 118.300 167.700 120.100 167.900 ;
        RECT 118.600 167.200 119.000 167.400 ;
        RECT 120.600 167.200 120.900 167.900 ;
        RECT 121.400 167.800 121.800 168.600 ;
        RECT 122.300 167.200 122.600 168.900 ;
        RECT 123.800 167.800 124.200 168.600 ;
        RECT 124.700 167.200 125.000 168.900 ;
        RECT 126.200 167.900 126.600 169.900 ;
        RECT 127.000 168.000 127.400 169.900 ;
        RECT 128.600 168.000 129.000 169.900 ;
        RECT 127.000 167.900 129.000 168.000 ;
        RECT 129.400 167.900 129.800 169.900 ;
        RECT 131.600 168.100 132.400 169.900 ;
        RECT 126.300 167.200 126.600 167.900 ;
        RECT 127.100 167.700 128.900 167.900 ;
        RECT 129.400 167.600 130.500 167.900 ;
        RECT 131.000 167.700 131.800 167.800 ;
        RECT 130.100 167.500 130.500 167.600 ;
        RECT 130.800 167.400 131.800 167.700 ;
        RECT 128.200 167.200 128.600 167.400 ;
        RECT 130.800 167.200 131.100 167.400 ;
        RECT 116.800 166.900 117.700 167.100 ;
        RECT 116.900 166.800 117.700 166.900 ;
        RECT 118.200 166.900 119.000 167.200 ;
        RECT 118.200 166.800 118.600 166.900 ;
        RECT 119.700 166.800 121.000 167.200 ;
        RECT 122.200 166.800 122.600 167.200 ;
        RECT 124.600 166.800 125.000 167.200 ;
        RECT 126.200 166.800 127.500 167.200 ;
        RECT 128.200 166.900 129.000 167.200 ;
        RECT 128.600 166.800 129.000 166.900 ;
        RECT 129.400 166.900 131.100 167.200 ;
        RECT 129.400 166.800 130.200 166.900 ;
        RECT 115.800 165.800 116.600 166.200 ;
        RECT 115.000 164.800 115.400 165.600 ;
        RECT 117.400 165.200 117.700 166.800 ;
        RECT 119.000 165.800 119.400 166.600 ;
        RECT 119.700 166.100 120.000 166.800 ;
        RECT 121.400 166.100 121.800 166.200 ;
        RECT 119.700 165.800 121.800 166.100 ;
        RECT 117.400 164.800 117.800 165.200 ;
        RECT 119.700 165.100 120.000 165.800 ;
        RECT 120.600 165.100 121.000 165.200 ;
        RECT 122.300 165.100 122.600 166.800 ;
        RECT 123.000 166.100 123.400 166.200 ;
        RECT 123.800 166.100 124.200 166.200 ;
        RECT 123.000 165.800 124.200 166.100 ;
        RECT 123.000 165.400 123.400 165.800 ;
        RECT 124.700 165.200 125.000 166.800 ;
        RECT 125.400 165.400 125.800 166.200 ;
        RECT 124.600 165.100 125.000 165.200 ;
        RECT 126.200 165.100 126.600 165.200 ;
        RECT 127.200 165.100 127.500 166.800 ;
        RECT 131.400 166.700 131.800 167.100 ;
        RECT 127.800 166.100 128.200 166.600 ;
        RECT 131.400 166.400 131.700 166.700 ;
        RECT 128.600 166.100 129.000 166.200 ;
        RECT 127.800 165.800 129.000 166.100 ;
        RECT 130.400 166.100 131.700 166.400 ;
        RECT 132.100 166.400 132.400 168.100 ;
        RECT 134.200 167.900 134.600 169.900 ;
        RECT 135.800 168.000 136.200 169.900 ;
        RECT 132.700 167.400 133.100 167.800 ;
        RECT 133.400 167.600 134.600 167.900 ;
        RECT 135.700 167.600 136.200 168.000 ;
        RECT 133.400 167.500 133.800 167.600 ;
        RECT 132.800 167.200 133.100 167.400 ;
        RECT 132.800 166.800 133.200 167.200 ;
        RECT 133.800 167.100 134.600 167.200 ;
        RECT 135.700 167.100 136.100 167.600 ;
        RECT 136.600 167.300 137.000 169.900 ;
        RECT 139.800 168.300 140.200 169.900 ;
        RECT 140.600 168.500 141.000 169.900 ;
        RECT 141.400 168.500 141.800 169.900 ;
        RECT 142.200 168.500 142.600 169.900 ;
        RECT 143.000 168.500 143.400 169.900 ;
        RECT 144.600 168.500 145.000 169.900 ;
        RECT 146.200 168.500 146.600 169.900 ;
        RECT 147.000 168.500 147.400 169.900 ;
        RECT 147.800 168.500 148.200 169.900 ;
        RECT 139.000 167.900 140.200 168.300 ;
        RECT 148.600 168.300 149.000 169.900 ;
        RECT 139.000 167.600 139.400 167.900 ;
        RECT 133.800 166.800 136.100 167.100 ;
        RECT 132.100 166.200 132.600 166.400 ;
        RECT 132.100 166.100 133.000 166.200 ;
        RECT 130.400 166.000 130.800 166.100 ;
        RECT 132.300 165.800 133.000 166.100 ;
        RECT 131.500 165.700 131.900 165.800 ;
        RECT 130.200 165.400 131.900 165.700 ;
        RECT 130.200 165.100 130.500 165.400 ;
        RECT 132.300 165.100 132.600 165.800 ;
        RECT 135.700 165.400 136.100 166.800 ;
        RECT 136.400 167.000 137.000 167.300 ;
        RECT 138.500 167.300 139.400 167.600 ;
        RECT 141.400 167.800 141.900 168.200 ;
        RECT 143.400 167.800 144.200 168.200 ;
        RECT 144.600 167.900 146.900 168.200 ;
        RECT 148.600 167.900 149.900 168.300 ;
        RECT 144.600 167.800 145.000 167.900 ;
        RECT 136.400 166.000 136.700 167.000 ;
        RECT 138.500 166.700 138.900 167.300 ;
        RECT 137.000 166.300 138.900 166.700 ;
        RECT 141.400 166.400 141.800 167.800 ;
        RECT 144.600 167.400 145.000 167.500 ;
        RECT 142.800 167.100 145.000 167.400 ;
        RECT 142.800 167.000 143.200 167.100 ;
        RECT 145.400 166.800 145.800 167.600 ;
        RECT 146.500 166.700 146.900 167.900 ;
        RECT 149.500 167.600 149.900 167.900 ;
        RECT 149.500 167.200 151.000 167.600 ;
        RECT 151.800 166.900 152.200 169.900 ;
        RECT 154.200 167.900 154.600 169.900 ;
        RECT 156.400 168.100 157.200 169.900 ;
        RECT 154.200 167.600 155.400 167.900 ;
        RECT 155.000 167.500 155.400 167.600 ;
        RECT 155.700 167.400 156.100 167.800 ;
        RECT 155.700 167.200 156.000 167.400 ;
        RECT 143.000 166.300 144.600 166.700 ;
        RECT 146.500 166.300 147.500 166.700 ;
        RECT 147.800 166.500 152.200 166.900 ;
        RECT 154.200 166.800 155.000 167.200 ;
        RECT 155.600 166.800 156.000 167.200 ;
        RECT 139.800 166.000 140.200 166.300 ;
        RECT 148.600 166.000 149.000 166.200 ;
        RECT 151.100 166.000 151.500 166.100 ;
        RECT 136.400 165.700 136.800 166.000 ;
        RECT 139.800 165.700 151.500 166.000 ;
        RECT 119.500 164.800 120.000 165.100 ;
        RECT 120.300 164.800 121.000 165.100 ;
        RECT 116.600 163.800 117.000 164.600 ;
        RECT 117.400 163.500 117.700 164.800 ;
        RECT 115.900 163.200 117.700 163.500 ;
        RECT 115.900 163.100 116.200 163.200 ;
        RECT 115.800 161.100 116.200 163.100 ;
        RECT 117.400 163.100 117.700 163.200 ;
        RECT 117.400 161.100 117.800 163.100 ;
        RECT 119.500 161.100 119.900 164.800 ;
        RECT 120.300 164.200 120.600 164.800 ;
        RECT 122.200 164.700 123.100 165.100 ;
        RECT 124.600 164.700 125.500 165.100 ;
        RECT 126.200 164.800 126.900 165.100 ;
        RECT 127.200 164.800 127.700 165.100 ;
        RECT 120.200 163.800 120.600 164.200 ;
        RECT 122.700 162.200 123.100 164.700 ;
        RECT 122.700 161.800 123.400 162.200 ;
        RECT 122.700 161.100 123.100 161.800 ;
        RECT 125.100 161.100 125.500 164.700 ;
        RECT 126.600 164.200 126.900 164.800 ;
        RECT 126.600 163.800 127.000 164.200 ;
        RECT 127.300 161.100 127.700 164.800 ;
        RECT 129.400 164.800 130.500 165.100 ;
        RECT 129.400 161.100 129.800 164.800 ;
        RECT 130.100 164.700 130.500 164.800 ;
        RECT 131.600 164.800 132.600 165.100 ;
        RECT 133.400 164.800 134.600 165.100 ;
        RECT 135.700 165.000 136.200 165.400 ;
        RECT 131.600 161.100 132.400 164.800 ;
        RECT 133.400 164.700 133.800 164.800 ;
        RECT 134.200 161.100 134.600 164.800 ;
        RECT 135.800 161.100 136.200 165.000 ;
        RECT 136.500 164.800 136.800 165.700 ;
        RECT 136.500 164.500 141.000 164.800 ;
        RECT 136.500 163.700 136.800 164.500 ;
        RECT 140.600 164.400 141.000 164.500 ;
        RECT 142.200 164.500 146.500 164.800 ;
        RECT 142.200 164.400 142.600 164.500 ;
        RECT 138.100 163.800 139.400 164.200 ;
        RECT 136.500 163.400 137.800 163.700 ;
        RECT 137.400 161.100 137.800 163.400 ;
        RECT 139.000 161.100 139.400 163.800 ;
        RECT 139.700 163.400 141.800 163.800 ;
        RECT 140.600 161.100 141.000 162.500 ;
        RECT 141.400 161.100 141.800 162.500 ;
        RECT 142.200 161.100 142.600 162.500 ;
        RECT 143.000 161.100 143.400 164.200 ;
        RECT 144.600 163.800 145.900 164.200 ;
        RECT 146.200 164.100 146.500 164.500 ;
        RECT 147.000 164.700 147.400 164.800 ;
        RECT 147.000 164.500 149.700 164.700 ;
        RECT 147.000 164.400 150.100 164.500 ;
        RECT 149.400 164.100 150.100 164.400 ;
        RECT 146.200 163.800 149.100 164.100 ;
        RECT 150.600 164.000 151.400 164.400 ;
        RECT 150.600 163.800 150.900 164.000 ;
        RECT 144.600 161.100 145.000 163.500 ;
        RECT 146.200 161.100 146.600 163.500 ;
        RECT 148.800 163.400 150.900 163.800 ;
        RECT 151.800 163.700 152.200 166.500 ;
        RECT 156.400 166.400 156.700 168.100 ;
        RECT 159.000 167.900 159.400 169.900 ;
        RECT 157.000 167.700 157.800 167.800 ;
        RECT 157.000 167.400 158.000 167.700 ;
        RECT 158.300 167.600 159.400 167.900 ;
        RECT 159.800 167.900 160.200 169.900 ;
        RECT 162.000 168.100 162.800 169.900 ;
        RECT 159.800 167.600 160.900 167.900 ;
        RECT 161.400 167.700 162.200 167.800 ;
        RECT 158.300 167.500 158.700 167.600 ;
        RECT 160.500 167.500 160.900 167.600 ;
        RECT 157.700 167.200 158.000 167.400 ;
        RECT 161.200 167.400 162.200 167.700 ;
        RECT 161.200 167.200 161.500 167.400 ;
        RECT 157.000 166.700 157.400 167.100 ;
        RECT 157.700 166.900 159.400 167.200 ;
        RECT 158.600 166.800 159.400 166.900 ;
        RECT 159.800 166.900 161.500 167.200 ;
        RECT 159.800 166.800 160.600 166.900 ;
        RECT 156.200 166.200 156.700 166.400 ;
        RECT 155.800 166.100 156.700 166.200 ;
        RECT 157.100 166.400 157.400 166.700 ;
        RECT 161.800 166.700 162.200 167.100 ;
        RECT 161.800 166.400 162.100 166.700 ;
        RECT 157.100 166.100 158.400 166.400 ;
        RECT 155.800 165.800 156.500 166.100 ;
        RECT 158.000 166.000 158.400 166.100 ;
        RECT 160.800 166.100 162.100 166.400 ;
        RECT 162.500 166.400 162.800 168.100 ;
        RECT 164.600 167.900 165.000 169.900 ;
        RECT 163.100 167.400 163.500 167.800 ;
        RECT 163.800 167.600 165.000 167.900 ;
        RECT 163.800 167.500 164.200 167.600 ;
        RECT 163.200 167.200 163.500 167.400 ;
        RECT 163.200 166.800 163.600 167.200 ;
        RECT 164.200 166.800 165.000 167.200 ;
        RECT 165.400 166.900 165.800 169.900 ;
        RECT 168.600 168.300 169.000 169.900 ;
        RECT 169.400 168.500 169.800 169.900 ;
        RECT 170.200 168.500 170.600 169.900 ;
        RECT 171.000 168.500 171.400 169.900 ;
        RECT 172.600 168.500 173.000 169.900 ;
        RECT 174.200 168.500 174.600 169.900 ;
        RECT 175.000 168.500 175.400 169.900 ;
        RECT 175.800 168.500 176.200 169.900 ;
        RECT 176.600 168.500 177.000 169.900 ;
        RECT 167.700 167.900 169.000 168.300 ;
        RECT 177.400 168.300 177.800 169.900 ;
        RECT 170.700 167.900 173.000 168.200 ;
        RECT 167.700 167.600 168.100 167.900 ;
        RECT 166.600 167.200 168.100 167.600 ;
        RECT 165.400 166.500 169.800 166.900 ;
        RECT 170.700 166.700 171.100 167.900 ;
        RECT 172.600 167.800 173.000 167.900 ;
        RECT 173.400 167.800 174.200 168.200 ;
        RECT 175.700 167.800 176.200 168.200 ;
        RECT 177.400 167.900 178.600 168.300 ;
        RECT 171.800 166.800 172.200 167.600 ;
        RECT 172.600 167.400 173.000 167.500 ;
        RECT 172.600 167.100 174.800 167.400 ;
        RECT 174.400 167.000 174.800 167.100 ;
        RECT 162.500 166.200 163.000 166.400 ;
        RECT 162.500 166.100 163.400 166.200 ;
        RECT 160.800 166.000 161.200 166.100 ;
        RECT 162.700 165.800 163.400 166.100 ;
        RECT 156.200 165.100 156.500 165.800 ;
        RECT 156.900 165.700 157.300 165.800 ;
        RECT 161.900 165.700 162.300 165.800 ;
        RECT 156.900 165.400 158.600 165.700 ;
        RECT 158.300 165.100 158.600 165.400 ;
        RECT 160.600 165.400 162.300 165.700 ;
        RECT 160.600 165.100 160.900 165.400 ;
        RECT 162.700 165.100 163.000 165.800 ;
        RECT 151.200 163.400 152.200 163.700 ;
        RECT 154.200 164.800 155.400 165.100 ;
        RECT 156.200 164.800 157.200 165.100 ;
        RECT 147.000 161.100 147.400 162.500 ;
        RECT 147.800 161.100 148.200 162.500 ;
        RECT 149.400 161.100 149.800 163.400 ;
        RECT 151.200 163.100 151.500 163.400 ;
        RECT 151.000 162.800 151.500 163.100 ;
        RECT 151.000 161.100 151.400 162.800 ;
        RECT 154.200 161.100 154.600 164.800 ;
        RECT 155.000 164.700 155.400 164.800 ;
        RECT 156.400 161.100 157.200 164.800 ;
        RECT 158.300 164.800 159.400 165.100 ;
        RECT 158.300 164.700 158.700 164.800 ;
        RECT 159.000 161.100 159.400 164.800 ;
        RECT 159.800 164.800 160.900 165.100 ;
        RECT 159.800 161.100 160.200 164.800 ;
        RECT 160.500 164.700 160.900 164.800 ;
        RECT 162.000 164.800 163.000 165.100 ;
        RECT 163.800 164.800 165.000 165.100 ;
        RECT 162.000 164.200 162.800 164.800 ;
        RECT 163.800 164.700 164.200 164.800 ;
        RECT 161.400 163.800 162.800 164.200 ;
        RECT 162.000 161.100 162.800 163.800 ;
        RECT 164.600 161.100 165.000 164.800 ;
        RECT 165.400 163.700 165.800 166.500 ;
        RECT 170.100 166.300 171.100 166.700 ;
        RECT 173.000 166.300 174.600 166.700 ;
        RECT 175.800 166.400 176.200 167.800 ;
        RECT 178.200 167.600 178.600 167.900 ;
        RECT 178.200 167.300 179.100 167.600 ;
        RECT 178.700 166.700 179.100 167.300 ;
        RECT 180.600 167.300 181.000 169.900 ;
        RECT 181.400 168.000 181.800 169.900 ;
        RECT 184.300 168.200 184.700 169.900 ;
        RECT 181.400 167.600 181.900 168.000 ;
        RECT 183.800 167.900 184.700 168.200 ;
        RECT 185.400 167.900 185.800 169.900 ;
        RECT 186.200 168.000 186.600 169.900 ;
        RECT 187.800 168.000 188.200 169.900 ;
        RECT 186.200 167.900 188.200 168.000 ;
        RECT 180.600 167.000 181.200 167.300 ;
        RECT 178.700 166.300 180.600 166.700 ;
        RECT 166.100 166.000 166.500 166.100 ;
        RECT 167.000 166.000 167.400 166.200 ;
        RECT 168.600 166.000 169.000 166.200 ;
        RECT 177.400 166.000 177.800 166.300 ;
        RECT 180.900 166.000 181.200 167.000 ;
        RECT 166.100 165.700 177.800 166.000 ;
        RECT 180.800 165.700 181.200 166.000 ;
        RECT 180.800 164.800 181.100 165.700 ;
        RECT 181.500 165.400 181.900 167.600 ;
        RECT 183.000 166.800 183.400 167.600 ;
        RECT 170.200 164.700 170.600 164.800 ;
        RECT 167.900 164.500 170.600 164.700 ;
        RECT 167.500 164.400 170.600 164.500 ;
        RECT 171.100 164.500 175.400 164.800 ;
        RECT 166.200 164.000 167.000 164.400 ;
        RECT 167.500 164.100 168.200 164.400 ;
        RECT 171.100 164.100 171.400 164.500 ;
        RECT 175.000 164.400 175.400 164.500 ;
        RECT 176.600 164.500 181.100 164.800 ;
        RECT 176.600 164.400 177.000 164.500 ;
        RECT 166.700 163.800 167.000 164.000 ;
        RECT 168.500 163.800 171.400 164.100 ;
        RECT 171.700 163.800 173.000 164.200 ;
        RECT 165.400 163.400 166.400 163.700 ;
        RECT 166.700 163.400 168.800 163.800 ;
        RECT 166.100 163.100 166.400 163.400 ;
        RECT 166.100 162.800 166.600 163.100 ;
        RECT 166.200 161.100 166.600 162.800 ;
        RECT 167.800 161.100 168.200 163.400 ;
        RECT 169.400 161.100 169.800 162.500 ;
        RECT 170.200 161.100 170.600 162.500 ;
        RECT 171.000 161.100 171.400 163.500 ;
        RECT 172.600 161.100 173.000 163.500 ;
        RECT 174.200 161.100 174.600 164.200 ;
        RECT 178.200 163.800 179.500 164.200 ;
        RECT 175.800 163.400 177.900 163.800 ;
        RECT 175.000 161.100 175.400 162.500 ;
        RECT 175.800 161.100 176.200 162.500 ;
        RECT 176.600 161.100 177.000 162.500 ;
        RECT 178.200 161.100 178.600 163.800 ;
        RECT 180.800 163.700 181.100 164.500 ;
        RECT 179.800 163.400 181.100 163.700 ;
        RECT 181.400 165.000 181.900 165.400 ;
        RECT 183.800 166.100 184.200 167.900 ;
        RECT 185.500 167.200 185.800 167.900 ;
        RECT 186.300 167.700 188.100 167.900 ;
        RECT 190.200 167.800 190.600 169.900 ;
        RECT 190.900 168.200 191.300 168.600 ;
        RECT 191.000 167.800 191.400 168.200 ;
        RECT 191.800 167.900 192.200 169.900 ;
        RECT 194.000 168.100 194.800 169.900 ;
        RECT 187.400 167.200 187.800 167.400 ;
        RECT 185.400 166.800 186.700 167.200 ;
        RECT 187.400 166.900 188.200 167.200 ;
        RECT 187.800 166.800 188.200 166.900 ;
        RECT 183.800 165.800 185.700 166.100 ;
        RECT 179.800 161.100 180.200 163.400 ;
        RECT 181.400 161.100 181.800 165.000 ;
        RECT 183.800 161.100 184.200 165.800 ;
        RECT 185.400 165.200 185.700 165.800 ;
        RECT 184.600 164.400 185.000 165.200 ;
        RECT 185.400 165.100 185.800 165.200 ;
        RECT 186.400 165.100 186.700 166.800 ;
        RECT 187.000 165.800 187.400 166.600 ;
        RECT 189.400 166.400 189.800 167.200 ;
        RECT 188.600 166.100 189.000 166.200 ;
        RECT 190.200 166.100 190.500 167.800 ;
        RECT 191.800 167.600 193.100 167.900 ;
        RECT 192.700 167.500 193.100 167.600 ;
        RECT 193.400 167.400 194.200 167.800 ;
        RECT 191.800 167.100 192.600 167.200 ;
        RECT 194.500 167.100 194.800 168.100 ;
        RECT 196.600 167.900 197.000 169.900 ;
        RECT 197.400 168.000 197.800 169.900 ;
        RECT 199.000 168.000 199.400 169.900 ;
        RECT 197.400 167.900 199.400 168.000 ;
        RECT 199.800 167.900 200.200 169.900 ;
        RECT 195.100 167.400 195.500 167.800 ;
        RECT 195.800 167.600 197.000 167.900 ;
        RECT 197.500 167.700 199.300 167.900 ;
        RECT 195.800 167.500 196.200 167.600 ;
        RECT 191.800 167.000 192.900 167.100 ;
        RECT 191.800 166.800 194.000 167.000 ;
        RECT 192.600 166.700 194.000 166.800 ;
        RECT 193.600 166.600 194.000 166.700 ;
        RECT 194.300 166.800 194.800 167.100 ;
        RECT 195.200 167.200 195.500 167.400 ;
        RECT 197.800 167.200 198.200 167.400 ;
        RECT 199.800 167.200 200.100 167.900 ;
        RECT 195.200 166.800 195.600 167.200 ;
        RECT 196.200 166.800 197.000 167.200 ;
        RECT 197.400 166.900 198.200 167.200 ;
        RECT 197.400 166.800 197.800 166.900 ;
        RECT 198.900 166.800 200.200 167.200 ;
        RECT 202.400 167.100 202.800 169.900 ;
        RECT 202.400 166.900 203.300 167.100 ;
        RECT 202.500 166.800 203.300 166.900 ;
        RECT 194.300 166.200 194.600 166.800 ;
        RECT 191.000 166.100 191.400 166.200 ;
        RECT 188.600 165.800 189.400 166.100 ;
        RECT 190.200 165.800 191.400 166.100 ;
        RECT 192.900 166.100 193.300 166.200 ;
        RECT 192.900 165.800 193.700 166.100 ;
        RECT 194.200 165.800 194.600 166.200 ;
        RECT 198.200 165.800 198.600 166.600 ;
        RECT 198.900 166.100 199.200 166.800 ;
        RECT 199.800 166.100 200.200 166.200 ;
        RECT 198.900 165.800 200.200 166.100 ;
        RECT 201.400 165.800 202.200 166.200 ;
        RECT 189.000 165.600 189.400 165.800 ;
        RECT 191.000 165.100 191.300 165.800 ;
        RECT 193.300 165.700 193.700 165.800 ;
        RECT 194.300 165.100 194.600 165.800 ;
        RECT 198.900 165.100 199.200 165.800 ;
        RECT 203.000 165.200 203.300 166.800 ;
        RECT 199.800 165.100 200.200 165.200 ;
        RECT 185.400 164.800 186.100 165.100 ;
        RECT 186.400 164.800 186.900 165.100 ;
        RECT 185.800 164.200 186.100 164.800 ;
        RECT 185.800 163.800 186.200 164.200 ;
        RECT 186.500 161.100 186.900 164.800 ;
        RECT 188.600 164.800 190.600 165.100 ;
        RECT 188.600 161.100 189.000 164.800 ;
        RECT 190.200 161.100 190.600 164.800 ;
        RECT 191.000 161.100 191.400 165.100 ;
        RECT 191.800 164.800 193.100 165.100 ;
        RECT 191.800 161.100 192.200 164.800 ;
        RECT 192.700 164.700 193.100 164.800 ;
        RECT 194.000 161.100 194.800 165.100 ;
        RECT 195.800 164.800 197.000 165.100 ;
        RECT 195.800 164.700 196.200 164.800 ;
        RECT 196.600 161.100 197.000 164.800 ;
        RECT 198.700 164.800 199.200 165.100 ;
        RECT 199.500 164.800 200.200 165.100 ;
        RECT 203.000 164.800 203.400 165.200 ;
        RECT 198.700 161.100 199.100 164.800 ;
        RECT 199.500 164.200 199.800 164.800 ;
        RECT 199.400 164.100 199.800 164.200 ;
        RECT 199.400 163.800 201.700 164.100 ;
        RECT 202.200 163.800 202.600 164.600 ;
        RECT 201.400 163.500 201.700 163.800 ;
        RECT 203.000 163.500 203.300 164.800 ;
        RECT 201.400 163.200 203.300 163.500 ;
        RECT 201.400 161.100 201.800 163.200 ;
        RECT 203.000 163.100 203.300 163.200 ;
        RECT 203.000 161.100 203.400 163.100 ;
        RECT 203.800 161.100 204.200 169.900 ;
        RECT 204.600 167.800 205.000 168.600 ;
        RECT 2.200 156.200 2.600 159.900 ;
        RECT 4.600 156.200 5.000 159.900 ;
        RECT 1.500 155.900 2.600 156.200 ;
        RECT 3.900 155.900 5.000 156.200 ;
        RECT 1.500 155.600 1.800 155.900 ;
        RECT 3.900 155.600 4.200 155.900 ;
        RECT 1.200 155.200 1.800 155.600 ;
        RECT 3.600 155.200 4.200 155.600 ;
        RECT 5.400 155.700 5.800 159.900 ;
        RECT 7.600 158.200 8.000 159.900 ;
        RECT 7.000 157.900 8.000 158.200 ;
        RECT 9.800 157.900 10.200 159.900 ;
        RECT 11.900 157.900 12.500 159.900 ;
        RECT 7.000 157.500 7.400 157.900 ;
        RECT 9.800 157.600 10.100 157.900 ;
        RECT 8.700 157.300 10.500 157.600 ;
        RECT 11.800 157.500 12.200 157.900 ;
        RECT 8.700 157.200 9.100 157.300 ;
        RECT 10.100 157.200 10.500 157.300 ;
        RECT 7.000 156.500 7.400 156.600 ;
        RECT 9.300 156.500 9.700 156.600 ;
        RECT 7.000 156.200 9.700 156.500 ;
        RECT 10.000 156.500 11.100 156.800 ;
        RECT 10.000 155.900 10.300 156.500 ;
        RECT 10.700 156.400 11.100 156.500 ;
        RECT 11.900 156.600 12.600 157.000 ;
        RECT 11.900 156.100 12.200 156.600 ;
        RECT 7.900 155.700 10.300 155.900 ;
        RECT 5.400 155.600 10.300 155.700 ;
        RECT 11.000 155.800 12.200 156.100 ;
        RECT 5.400 155.500 8.300 155.600 ;
        RECT 5.400 155.400 8.200 155.500 ;
        RECT 1.500 153.700 1.800 155.200 ;
        RECT 2.200 154.400 2.600 155.200 ;
        RECT 3.900 153.700 4.200 155.200 ;
        RECT 4.600 154.400 5.000 155.200 ;
        RECT 8.600 155.100 9.000 155.200 ;
        RECT 10.200 155.100 10.600 155.200 ;
        RECT 6.500 154.800 10.600 155.100 ;
        RECT 6.500 154.700 6.900 154.800 ;
        RECT 7.300 154.200 7.700 154.300 ;
        RECT 11.000 154.200 11.300 155.800 ;
        RECT 14.200 155.600 14.600 159.900 ;
        RECT 16.300 156.300 16.700 159.900 ;
        RECT 15.800 155.900 16.700 156.300 ;
        RECT 18.200 156.000 18.600 159.900 ;
        RECT 19.800 157.600 20.200 159.900 ;
        RECT 12.500 155.300 14.600 155.600 ;
        RECT 12.500 155.200 12.900 155.300 ;
        RECT 13.300 154.900 13.700 155.000 ;
        RECT 11.800 154.600 13.700 154.900 ;
        RECT 11.800 154.500 12.200 154.600 ;
        RECT 5.800 153.900 11.300 154.200 ;
        RECT 5.800 153.800 6.600 153.900 ;
        RECT 1.500 153.400 2.600 153.700 ;
        RECT 3.900 153.400 5.000 153.700 ;
        RECT 2.200 151.100 2.600 153.400 ;
        RECT 4.600 151.100 5.000 153.400 ;
        RECT 5.400 151.100 5.800 153.500 ;
        RECT 7.900 152.800 8.200 153.900 ;
        RECT 9.400 153.800 9.800 153.900 ;
        RECT 10.700 153.800 11.100 153.900 ;
        RECT 14.200 153.600 14.600 155.300 ;
        RECT 15.900 154.200 16.200 155.900 ;
        RECT 18.100 155.600 18.600 156.000 ;
        RECT 18.900 157.300 20.200 157.600 ;
        RECT 18.900 156.500 19.200 157.300 ;
        RECT 21.400 157.200 21.800 159.900 ;
        RECT 23.000 158.500 23.400 159.900 ;
        RECT 23.800 158.500 24.200 159.900 ;
        RECT 24.600 158.500 25.000 159.900 ;
        RECT 22.100 157.200 24.200 157.600 ;
        RECT 20.500 156.800 21.800 157.200 ;
        RECT 25.400 156.800 25.800 159.900 ;
        RECT 27.000 157.500 27.400 159.900 ;
        RECT 28.600 157.500 29.000 159.900 ;
        RECT 29.400 158.500 29.800 159.900 ;
        RECT 30.200 158.500 30.600 159.900 ;
        RECT 31.800 157.600 32.200 159.900 ;
        RECT 33.400 158.200 33.800 159.900 ;
        RECT 33.400 157.900 33.900 158.200 ;
        RECT 33.600 157.600 33.900 157.900 ;
        RECT 31.200 157.200 33.300 157.600 ;
        RECT 33.600 157.300 34.600 157.600 ;
        RECT 27.000 156.800 28.300 157.200 ;
        RECT 28.600 156.900 31.500 157.200 ;
        RECT 33.000 157.000 33.300 157.200 ;
        RECT 23.000 156.500 23.400 156.600 ;
        RECT 18.900 156.200 23.400 156.500 ;
        RECT 24.600 156.500 25.000 156.600 ;
        RECT 28.600 156.500 28.900 156.900 ;
        RECT 31.800 156.600 32.500 156.900 ;
        RECT 33.000 156.600 33.800 157.000 ;
        RECT 24.600 156.200 28.900 156.500 ;
        RECT 29.400 156.500 32.500 156.600 ;
        RECT 29.400 156.300 32.100 156.500 ;
        RECT 29.400 156.200 29.800 156.300 ;
        RECT 16.600 154.800 17.000 155.600 ;
        RECT 15.800 153.800 16.200 154.200 ;
        RECT 12.700 153.300 14.600 153.600 ;
        RECT 12.700 153.200 13.100 153.300 ;
        RECT 14.200 153.100 14.600 153.300 ;
        RECT 15.000 153.100 15.400 153.200 ;
        RECT 14.200 152.800 15.400 153.100 ;
        RECT 7.000 152.100 7.400 152.500 ;
        RECT 7.800 152.400 8.200 152.800 ;
        RECT 8.700 152.700 9.100 152.800 ;
        RECT 8.700 152.400 10.100 152.700 ;
        RECT 9.800 152.100 10.100 152.400 ;
        RECT 11.800 152.100 12.200 152.500 ;
        RECT 7.000 151.800 8.000 152.100 ;
        RECT 7.600 151.100 8.000 151.800 ;
        RECT 9.800 151.100 10.200 152.100 ;
        RECT 11.800 151.800 12.500 152.100 ;
        RECT 11.900 151.100 12.500 151.800 ;
        RECT 14.200 151.100 14.600 152.800 ;
        RECT 15.000 152.400 15.400 152.800 ;
        RECT 15.900 152.200 16.200 153.800 ;
        RECT 18.100 153.400 18.500 155.600 ;
        RECT 18.900 155.300 19.200 156.200 ;
        RECT 18.800 155.000 19.200 155.300 ;
        RECT 22.200 155.000 33.900 155.300 ;
        RECT 18.800 154.000 19.100 155.000 ;
        RECT 22.200 154.700 22.600 155.000 ;
        RECT 31.000 154.800 31.400 155.000 ;
        RECT 33.400 154.900 33.900 155.000 ;
        RECT 33.400 154.800 33.800 154.900 ;
        RECT 19.400 154.300 21.300 154.700 ;
        RECT 18.800 153.700 19.400 154.000 ;
        RECT 18.100 153.000 18.600 153.400 ;
        RECT 15.800 151.100 16.200 152.200 ;
        RECT 18.200 151.100 18.600 153.000 ;
        RECT 19.000 151.100 19.400 153.700 ;
        RECT 20.900 153.700 21.300 154.300 ;
        RECT 20.900 153.400 21.800 153.700 ;
        RECT 21.400 153.100 21.800 153.400 ;
        RECT 23.800 153.200 24.200 154.600 ;
        RECT 25.400 154.300 27.000 154.700 ;
        RECT 28.900 154.300 29.900 154.700 ;
        RECT 34.200 154.500 34.600 157.300 ;
        RECT 35.000 156.200 35.400 159.900 ;
        RECT 36.600 156.200 37.000 159.900 ;
        RECT 35.000 155.900 37.000 156.200 ;
        RECT 37.400 155.900 37.800 159.900 ;
        RECT 38.500 156.300 38.900 159.900 ;
        RECT 38.500 155.900 39.400 156.300 ;
        RECT 35.400 155.200 35.800 155.400 ;
        RECT 37.400 155.200 37.700 155.900 ;
        RECT 35.000 154.900 35.800 155.200 ;
        RECT 36.600 154.900 37.800 155.200 ;
        RECT 35.000 154.800 35.400 154.900 ;
        RECT 25.200 153.900 25.600 154.000 ;
        RECT 25.200 153.600 27.400 153.900 ;
        RECT 27.000 153.500 27.400 153.600 ;
        RECT 27.800 153.400 28.200 154.200 ;
        RECT 21.400 152.700 22.600 153.100 ;
        RECT 23.800 152.800 24.300 153.200 ;
        RECT 25.800 152.800 26.600 153.200 ;
        RECT 27.000 153.100 27.400 153.200 ;
        RECT 28.900 153.100 29.300 154.300 ;
        RECT 30.200 154.100 34.600 154.500 ;
        RECT 31.900 153.400 33.400 153.800 ;
        RECT 31.900 153.100 32.300 153.400 ;
        RECT 27.000 152.800 29.300 153.100 ;
        RECT 22.200 151.100 22.600 152.700 ;
        RECT 31.000 152.700 32.300 153.100 ;
        RECT 23.000 151.100 23.400 152.500 ;
        RECT 23.800 151.100 24.200 152.500 ;
        RECT 24.600 151.100 25.000 152.500 ;
        RECT 25.400 151.100 25.800 152.500 ;
        RECT 27.000 151.100 27.400 152.500 ;
        RECT 28.600 151.100 29.000 152.500 ;
        RECT 29.400 151.100 29.800 152.500 ;
        RECT 30.200 151.100 30.600 152.500 ;
        RECT 31.000 151.100 31.400 152.700 ;
        RECT 34.200 151.100 34.600 154.100 ;
        RECT 35.800 153.800 36.200 154.600 ;
        RECT 36.600 153.100 36.900 154.900 ;
        RECT 37.400 154.800 37.800 154.900 ;
        RECT 38.200 154.800 38.600 155.600 ;
        RECT 39.000 154.200 39.300 155.900 ;
        RECT 40.600 155.700 41.000 159.900 ;
        RECT 42.800 158.200 43.200 159.900 ;
        RECT 42.200 157.900 43.200 158.200 ;
        RECT 45.000 157.900 45.400 159.900 ;
        RECT 47.100 157.900 47.700 159.900 ;
        RECT 42.200 157.500 42.600 157.900 ;
        RECT 45.000 157.600 45.300 157.900 ;
        RECT 43.900 157.300 45.700 157.600 ;
        RECT 47.000 157.500 47.400 157.900 ;
        RECT 43.900 157.200 44.300 157.300 ;
        RECT 45.300 157.200 45.700 157.300 ;
        RECT 42.200 156.500 42.600 156.600 ;
        RECT 44.500 156.500 44.900 156.600 ;
        RECT 42.200 156.200 44.900 156.500 ;
        RECT 45.200 156.500 46.300 156.800 ;
        RECT 45.200 155.900 45.500 156.500 ;
        RECT 45.900 156.400 46.300 156.500 ;
        RECT 47.100 156.600 47.800 157.000 ;
        RECT 47.100 156.100 47.400 156.600 ;
        RECT 43.100 155.700 45.500 155.900 ;
        RECT 40.600 155.600 45.500 155.700 ;
        RECT 46.200 155.800 47.400 156.100 ;
        RECT 40.600 155.500 43.500 155.600 ;
        RECT 40.600 155.400 43.400 155.500 ;
        RECT 43.800 155.100 44.200 155.200 ;
        RECT 41.700 154.800 44.200 155.100 ;
        RECT 41.700 154.700 42.100 154.800 ;
        RECT 42.500 154.200 42.900 154.300 ;
        RECT 46.200 154.200 46.500 155.800 ;
        RECT 49.400 155.600 49.800 159.900 ;
        RECT 53.100 156.200 53.500 159.900 ;
        RECT 53.800 156.800 54.200 157.200 ;
        RECT 53.900 156.200 54.200 156.800 ;
        RECT 52.600 155.800 53.600 156.200 ;
        RECT 53.900 156.100 54.600 156.200 ;
        RECT 55.800 156.100 56.200 159.900 ;
        RECT 53.900 155.900 56.200 156.100 ;
        RECT 54.200 155.800 56.200 155.900 ;
        RECT 56.600 155.800 57.000 156.600 ;
        RECT 57.400 156.200 57.800 159.900 ;
        RECT 59.000 156.200 59.400 159.900 ;
        RECT 57.400 155.900 59.400 156.200 ;
        RECT 59.800 155.900 60.200 159.900 ;
        RECT 47.700 155.300 49.800 155.600 ;
        RECT 47.700 155.200 48.100 155.300 ;
        RECT 48.500 154.900 48.900 155.000 ;
        RECT 47.000 154.600 48.900 154.900 ;
        RECT 47.000 154.500 47.400 154.600 ;
        RECT 39.000 153.800 39.400 154.200 ;
        RECT 41.000 153.900 46.500 154.200 ;
        RECT 41.000 153.800 41.800 153.900 ;
        RECT 37.400 153.100 37.800 153.200 ;
        RECT 39.000 153.100 39.300 153.800 ;
        RECT 36.600 151.100 37.000 153.100 ;
        RECT 37.400 152.800 39.300 153.100 ;
        RECT 37.300 152.400 37.700 152.800 ;
        RECT 39.000 152.100 39.300 152.800 ;
        RECT 39.800 152.400 40.200 153.200 ;
        RECT 39.000 151.100 39.400 152.100 ;
        RECT 40.600 151.100 41.000 153.500 ;
        RECT 43.100 152.800 43.400 153.900 ;
        RECT 44.600 153.800 45.000 153.900 ;
        RECT 45.900 153.800 46.300 153.900 ;
        RECT 49.400 153.600 49.800 155.300 ;
        RECT 51.800 155.100 52.200 155.200 ;
        RECT 52.600 155.100 53.000 155.200 ;
        RECT 51.800 154.800 53.000 155.100 ;
        RECT 52.600 154.400 53.000 154.800 ;
        RECT 53.300 154.200 53.600 155.800 ;
        RECT 51.800 154.100 52.200 154.200 ;
        RECT 51.800 153.800 52.600 154.100 ;
        RECT 53.300 153.800 54.600 154.200 ;
        RECT 52.200 153.600 52.600 153.800 ;
        RECT 47.900 153.300 49.800 153.600 ;
        RECT 47.900 153.200 48.300 153.300 ;
        RECT 42.200 152.100 42.600 152.500 ;
        RECT 43.000 152.400 43.400 152.800 ;
        RECT 43.900 152.700 44.300 152.800 ;
        RECT 43.900 152.400 45.300 152.700 ;
        RECT 45.000 152.100 45.300 152.400 ;
        RECT 47.000 152.100 47.400 152.500 ;
        RECT 42.200 151.800 43.200 152.100 ;
        RECT 42.800 151.100 43.200 151.800 ;
        RECT 45.000 151.100 45.400 152.100 ;
        RECT 47.000 151.800 47.700 152.100 ;
        RECT 47.100 151.100 47.700 151.800 ;
        RECT 49.400 151.100 49.800 153.300 ;
        RECT 51.900 153.100 53.700 153.300 ;
        RECT 54.200 153.100 54.500 153.800 ;
        RECT 55.000 153.400 55.400 154.200 ;
        RECT 55.800 153.100 56.200 155.800 ;
        RECT 57.800 155.200 58.200 155.400 ;
        RECT 59.800 155.200 60.100 155.900 ;
        RECT 60.600 155.700 61.000 159.900 ;
        RECT 62.800 158.200 63.200 159.900 ;
        RECT 62.200 157.900 63.200 158.200 ;
        RECT 65.000 157.900 65.400 159.900 ;
        RECT 67.100 157.900 67.700 159.900 ;
        RECT 62.200 157.500 62.600 157.900 ;
        RECT 65.000 157.600 65.300 157.900 ;
        RECT 63.900 157.300 65.700 157.600 ;
        RECT 67.000 157.500 67.400 157.900 ;
        RECT 63.900 157.200 64.300 157.300 ;
        RECT 65.300 157.200 65.700 157.300 ;
        RECT 62.200 156.500 62.600 156.600 ;
        RECT 64.500 156.500 64.900 156.600 ;
        RECT 62.200 156.200 64.900 156.500 ;
        RECT 65.200 156.500 66.300 156.800 ;
        RECT 65.200 155.900 65.500 156.500 ;
        RECT 65.900 156.400 66.300 156.500 ;
        RECT 67.100 156.600 67.800 157.000 ;
        RECT 67.100 156.100 67.400 156.600 ;
        RECT 63.100 155.700 65.500 155.900 ;
        RECT 60.600 155.600 65.500 155.700 ;
        RECT 66.200 155.800 67.400 156.100 ;
        RECT 60.600 155.500 63.500 155.600 ;
        RECT 60.600 155.400 63.400 155.500 ;
        RECT 66.200 155.200 66.500 155.800 ;
        RECT 69.400 155.600 69.800 159.900 ;
        RECT 71.500 156.200 71.900 159.900 ;
        RECT 72.200 156.800 72.600 157.200 ;
        RECT 72.300 156.200 72.600 156.800 ;
        RECT 71.500 155.900 72.000 156.200 ;
        RECT 72.300 155.900 73.000 156.200 ;
        RECT 67.700 155.300 69.800 155.600 ;
        RECT 67.700 155.200 68.100 155.300 ;
        RECT 57.400 154.900 58.200 155.200 ;
        RECT 59.000 154.900 60.200 155.200 ;
        RECT 63.800 155.100 64.200 155.200 ;
        RECT 57.400 154.800 57.800 154.900 ;
        RECT 58.200 153.800 58.600 154.600 ;
        RECT 59.000 153.100 59.300 154.900 ;
        RECT 59.800 154.800 60.200 154.900 ;
        RECT 61.700 154.800 64.200 155.100 ;
        RECT 66.200 154.800 66.600 155.200 ;
        RECT 68.500 154.900 68.900 155.000 ;
        RECT 59.800 154.200 60.100 154.800 ;
        RECT 61.700 154.700 62.100 154.800 ;
        RECT 63.000 154.700 63.400 154.800 ;
        RECT 62.500 154.200 62.900 154.300 ;
        RECT 66.200 154.200 66.500 154.800 ;
        RECT 67.000 154.600 68.900 154.900 ;
        RECT 67.000 154.500 67.400 154.600 ;
        RECT 59.800 153.800 60.200 154.200 ;
        RECT 61.000 153.900 66.500 154.200 ;
        RECT 61.000 153.800 61.800 153.900 ;
        RECT 51.800 153.000 53.800 153.100 ;
        RECT 51.800 151.100 52.200 153.000 ;
        RECT 53.400 151.100 53.800 153.000 ;
        RECT 54.200 151.100 54.600 153.100 ;
        RECT 55.800 152.800 56.700 153.100 ;
        RECT 56.300 151.100 56.700 152.800 ;
        RECT 59.000 151.100 59.400 153.100 ;
        RECT 59.800 152.800 60.200 153.200 ;
        RECT 59.700 152.400 60.100 152.800 ;
        RECT 60.600 151.100 61.000 153.500 ;
        RECT 63.100 152.800 63.400 153.900 ;
        RECT 65.900 153.800 66.300 153.900 ;
        RECT 69.400 153.600 69.800 155.300 ;
        RECT 71.700 155.200 72.000 155.900 ;
        RECT 72.600 155.800 73.000 155.900 ;
        RECT 73.400 155.800 73.800 156.600 ;
        RECT 71.000 154.400 71.400 155.200 ;
        RECT 71.700 154.800 72.200 155.200 ;
        RECT 72.600 155.100 72.900 155.800 ;
        RECT 74.200 155.100 74.600 159.900 ;
        RECT 72.600 154.800 74.600 155.100 ;
        RECT 71.700 154.200 72.000 154.800 ;
        RECT 70.200 154.100 70.600 154.200 ;
        RECT 70.200 153.800 71.000 154.100 ;
        RECT 71.700 153.800 73.000 154.200 ;
        RECT 70.600 153.600 71.000 153.800 ;
        RECT 67.900 153.300 69.800 153.600 ;
        RECT 67.900 153.200 68.300 153.300 ;
        RECT 62.200 152.100 62.600 152.500 ;
        RECT 63.000 152.400 63.400 152.800 ;
        RECT 63.900 152.700 64.300 152.800 ;
        RECT 63.900 152.400 65.300 152.700 ;
        RECT 65.000 152.100 65.300 152.400 ;
        RECT 67.000 152.100 67.400 152.500 ;
        RECT 62.200 151.800 63.200 152.100 ;
        RECT 62.800 151.100 63.200 151.800 ;
        RECT 65.000 151.100 65.400 152.100 ;
        RECT 67.000 151.800 67.700 152.100 ;
        RECT 67.100 151.100 67.700 151.800 ;
        RECT 69.400 151.100 69.800 153.300 ;
        RECT 70.300 153.100 72.100 153.300 ;
        RECT 72.600 153.100 72.900 153.800 ;
        RECT 74.200 153.100 74.600 154.800 ;
        RECT 75.000 153.400 75.400 154.200 ;
        RECT 75.800 153.400 76.200 154.200 ;
        RECT 70.200 153.000 72.200 153.100 ;
        RECT 70.200 151.100 70.600 153.000 ;
        RECT 71.800 151.100 72.200 153.000 ;
        RECT 72.600 151.100 73.000 153.100 ;
        RECT 73.700 152.800 74.600 153.100 ;
        RECT 76.600 153.100 77.000 159.900 ;
        RECT 79.000 158.200 79.400 159.900 ;
        RECT 78.900 157.900 79.400 158.200 ;
        RECT 78.900 157.600 79.200 157.900 ;
        RECT 80.600 157.600 81.000 159.900 ;
        RECT 82.200 158.500 82.600 159.900 ;
        RECT 83.000 158.500 83.400 159.900 ;
        RECT 78.200 157.300 79.200 157.600 ;
        RECT 77.400 155.800 77.800 156.600 ;
        RECT 78.200 154.500 78.600 157.300 ;
        RECT 79.500 157.200 81.600 157.600 ;
        RECT 83.800 157.500 84.200 159.900 ;
        RECT 85.400 157.500 85.800 159.900 ;
        RECT 79.500 157.000 79.800 157.200 ;
        RECT 79.000 156.600 79.800 157.000 ;
        RECT 81.300 156.900 84.200 157.200 ;
        RECT 80.300 156.600 81.000 156.900 ;
        RECT 80.300 156.500 83.400 156.600 ;
        RECT 80.700 156.300 83.400 156.500 ;
        RECT 83.000 156.200 83.400 156.300 ;
        RECT 83.900 156.500 84.200 156.900 ;
        RECT 84.500 156.800 85.800 157.200 ;
        RECT 87.000 156.800 87.400 159.900 ;
        RECT 87.800 158.500 88.200 159.900 ;
        RECT 88.600 158.500 89.000 159.900 ;
        RECT 89.400 158.500 89.800 159.900 ;
        RECT 88.600 157.200 90.700 157.600 ;
        RECT 91.000 157.200 91.400 159.900 ;
        RECT 92.600 157.600 93.000 159.900 ;
        RECT 92.600 157.300 93.900 157.600 ;
        RECT 91.000 156.800 92.300 157.200 ;
        RECT 87.800 156.500 88.200 156.600 ;
        RECT 83.900 156.200 88.200 156.500 ;
        RECT 89.400 156.500 89.800 156.600 ;
        RECT 93.600 156.500 93.900 157.300 ;
        RECT 89.400 156.200 93.900 156.500 ;
        RECT 93.600 155.300 93.900 156.200 ;
        RECT 94.200 156.100 94.600 159.900 ;
        RECT 96.900 157.200 97.300 159.900 ;
        RECT 96.200 156.800 96.600 157.200 ;
        RECT 96.900 156.800 97.800 157.200 ;
        RECT 96.200 156.200 96.500 156.800 ;
        RECT 96.900 156.200 97.300 156.800 ;
        RECT 95.800 156.100 96.500 156.200 ;
        RECT 94.200 155.900 96.500 156.100 ;
        RECT 96.800 155.900 97.300 156.200 ;
        RECT 99.300 156.300 99.700 159.900 ;
        RECT 99.300 155.900 100.200 156.300 ;
        RECT 94.200 155.800 96.200 155.900 ;
        RECT 94.200 155.600 94.700 155.800 ;
        RECT 78.900 155.000 90.600 155.300 ;
        RECT 93.600 155.000 94.000 155.300 ;
        RECT 78.900 154.900 79.300 155.000 ;
        RECT 81.400 154.800 81.800 155.000 ;
        RECT 90.200 154.700 90.600 155.000 ;
        RECT 78.200 154.100 82.600 154.500 ;
        RECT 82.900 154.300 83.900 154.700 ;
        RECT 85.800 154.300 87.400 154.700 ;
        RECT 76.600 152.800 77.500 153.100 ;
        RECT 73.700 151.100 74.100 152.800 ;
        RECT 77.100 151.100 77.500 152.800 ;
        RECT 78.200 151.100 78.600 154.100 ;
        RECT 79.400 153.400 80.900 153.800 ;
        RECT 80.500 153.100 80.900 153.400 ;
        RECT 83.500 153.100 83.900 154.300 ;
        RECT 84.600 153.400 85.000 154.200 ;
        RECT 87.200 153.900 87.600 154.000 ;
        RECT 85.400 153.600 87.600 153.900 ;
        RECT 85.400 153.500 85.800 153.600 ;
        RECT 88.600 153.200 89.000 154.600 ;
        RECT 91.500 154.300 93.400 154.700 ;
        RECT 91.500 153.700 91.900 154.300 ;
        RECT 93.700 154.000 94.000 155.000 ;
        RECT 85.400 153.100 85.800 153.200 ;
        RECT 80.500 152.700 81.800 153.100 ;
        RECT 83.500 152.800 85.800 153.100 ;
        RECT 86.200 152.800 87.000 153.200 ;
        RECT 88.500 152.800 89.000 153.200 ;
        RECT 91.000 153.400 91.900 153.700 ;
        RECT 93.400 153.700 94.000 154.000 ;
        RECT 91.000 153.100 91.400 153.400 ;
        RECT 81.400 151.100 81.800 152.700 ;
        RECT 90.200 152.700 91.400 153.100 ;
        RECT 82.200 151.100 82.600 152.500 ;
        RECT 83.000 151.100 83.400 152.500 ;
        RECT 83.800 151.100 84.200 152.500 ;
        RECT 85.400 151.100 85.800 152.500 ;
        RECT 87.000 151.100 87.400 152.500 ;
        RECT 87.800 151.100 88.200 152.500 ;
        RECT 88.600 151.100 89.000 152.500 ;
        RECT 89.400 151.100 89.800 152.500 ;
        RECT 90.200 151.100 90.600 152.700 ;
        RECT 93.400 151.100 93.800 153.700 ;
        RECT 94.300 153.400 94.700 155.600 ;
        RECT 96.800 154.200 97.100 155.900 ;
        RECT 97.400 155.100 97.800 155.200 ;
        RECT 99.000 155.100 99.400 155.600 ;
        RECT 97.400 154.800 99.400 155.100 ;
        RECT 97.400 154.400 97.800 154.800 ;
        RECT 99.800 154.200 100.100 155.900 ;
        RECT 95.800 153.800 97.100 154.200 ;
        RECT 98.200 154.100 98.600 154.200 ;
        RECT 97.800 153.800 98.600 154.100 ;
        RECT 99.800 153.800 100.200 154.200 ;
        RECT 94.200 153.000 94.700 153.400 ;
        RECT 95.900 153.100 96.200 153.800 ;
        RECT 97.800 153.600 98.200 153.800 ;
        RECT 96.700 153.100 98.500 153.300 ;
        RECT 94.200 151.100 94.600 153.000 ;
        RECT 95.800 151.100 96.200 153.100 ;
        RECT 96.600 153.000 98.600 153.100 ;
        RECT 96.600 151.100 97.000 153.000 ;
        RECT 98.200 151.100 98.600 153.000 ;
        RECT 99.800 152.200 100.100 153.800 ;
        RECT 100.600 153.100 101.000 153.200 ;
        RECT 103.000 153.100 103.400 153.200 ;
        RECT 100.600 152.800 103.400 153.100 ;
        RECT 100.600 152.400 101.000 152.800 ;
        RECT 103.000 152.400 103.400 152.800 ;
        RECT 99.800 151.100 100.200 152.200 ;
        RECT 103.800 151.100 104.200 159.900 ;
        RECT 105.900 156.300 106.300 159.900 ;
        RECT 105.400 155.900 106.300 156.300 ;
        RECT 105.500 154.200 105.800 155.900 ;
        RECT 106.200 154.800 106.600 155.600 ;
        RECT 105.400 154.100 105.800 154.200 ;
        RECT 107.000 154.100 107.400 154.200 ;
        RECT 105.400 153.800 107.400 154.100 ;
        RECT 104.600 152.400 105.000 153.200 ;
        RECT 105.500 152.100 105.800 153.800 ;
        RECT 107.000 153.400 107.400 153.800 ;
        RECT 107.800 153.100 108.200 159.900 ;
        RECT 108.600 155.800 109.000 156.600 ;
        RECT 110.700 156.300 111.100 159.900 ;
        RECT 110.200 155.900 111.100 156.300 ;
        RECT 111.800 156.200 112.200 159.900 ;
        RECT 113.400 156.400 113.800 159.900 ;
        RECT 111.800 155.900 113.100 156.200 ;
        RECT 113.400 155.900 113.900 156.400 ;
        RECT 110.300 154.200 110.600 155.900 ;
        RECT 111.000 154.800 111.400 155.600 ;
        RECT 111.800 154.800 112.300 155.200 ;
        RECT 111.900 154.400 112.300 154.800 ;
        RECT 112.800 154.900 113.100 155.900 ;
        RECT 112.800 154.500 113.300 154.900 ;
        RECT 110.200 153.800 110.600 154.200 ;
        RECT 110.300 153.200 110.600 153.800 ;
        RECT 112.800 153.700 113.100 154.500 ;
        RECT 113.600 154.200 113.900 155.900 ;
        RECT 113.400 153.800 113.900 154.200 ;
        RECT 109.400 153.100 109.800 153.200 ;
        RECT 107.800 152.800 109.800 153.100 ;
        RECT 110.200 152.800 110.600 153.200 ;
        RECT 105.400 151.100 105.800 152.100 ;
        RECT 108.300 151.100 108.700 152.800 ;
        RECT 109.400 152.400 109.800 152.800 ;
        RECT 110.300 152.100 110.600 152.800 ;
        RECT 110.200 151.100 110.600 152.100 ;
        RECT 111.800 153.400 113.100 153.700 ;
        RECT 111.800 151.100 112.200 153.400 ;
        RECT 113.600 153.200 113.900 153.800 ;
        RECT 115.000 154.800 115.400 155.200 ;
        RECT 115.000 154.200 115.300 154.800 ;
        RECT 115.000 153.400 115.400 154.200 ;
        RECT 113.400 152.800 113.900 153.200 ;
        RECT 115.800 153.100 116.200 159.900 ;
        RECT 116.600 155.800 117.000 156.600 ;
        RECT 118.700 156.300 119.100 159.900 ;
        RECT 118.200 155.900 119.100 156.300 ;
        RECT 118.300 154.200 118.600 155.900 ;
        RECT 119.000 154.800 119.400 155.600 ;
        RECT 118.200 153.800 118.600 154.200 ;
        RECT 117.400 153.100 117.800 153.200 ;
        RECT 115.800 152.800 117.800 153.100 ;
        RECT 113.400 151.100 113.800 152.800 ;
        RECT 116.300 151.100 116.700 152.800 ;
        RECT 117.400 152.400 117.800 152.800 ;
        RECT 118.300 152.200 118.600 153.800 ;
        RECT 119.800 153.400 120.200 154.200 ;
        RECT 120.600 153.100 121.000 159.900 ;
        RECT 121.400 155.800 121.800 156.600 ;
        RECT 122.200 153.400 122.600 154.200 ;
        RECT 123.000 153.100 123.400 159.900 ;
        RECT 123.800 156.100 124.200 156.600 ;
        RECT 124.600 156.100 125.000 156.200 ;
        RECT 123.800 155.800 125.000 156.100 ;
        RECT 125.400 156.000 125.800 159.900 ;
        RECT 127.000 157.600 127.400 159.900 ;
        RECT 125.300 155.600 125.800 156.000 ;
        RECT 126.100 157.300 127.400 157.600 ;
        RECT 126.100 156.500 126.400 157.300 ;
        RECT 128.600 157.200 129.000 159.900 ;
        RECT 130.200 158.500 130.600 159.900 ;
        RECT 131.000 158.500 131.400 159.900 ;
        RECT 131.800 158.500 132.200 159.900 ;
        RECT 129.300 157.200 131.400 157.600 ;
        RECT 127.700 156.800 129.000 157.200 ;
        RECT 132.600 156.800 133.000 159.900 ;
        RECT 134.200 157.500 134.600 159.900 ;
        RECT 135.800 157.500 136.200 159.900 ;
        RECT 136.600 158.500 137.000 159.900 ;
        RECT 137.400 158.500 137.800 159.900 ;
        RECT 139.000 157.600 139.400 159.900 ;
        RECT 140.600 158.200 141.000 159.900 ;
        RECT 140.600 157.900 141.100 158.200 ;
        RECT 140.800 157.600 141.100 157.900 ;
        RECT 138.400 157.200 140.500 157.600 ;
        RECT 140.800 157.300 141.800 157.600 ;
        RECT 134.200 156.800 135.500 157.200 ;
        RECT 135.800 156.900 138.700 157.200 ;
        RECT 140.200 157.000 140.500 157.200 ;
        RECT 130.200 156.500 130.600 156.600 ;
        RECT 126.100 156.200 130.600 156.500 ;
        RECT 131.800 156.500 132.200 156.600 ;
        RECT 135.800 156.500 136.100 156.900 ;
        RECT 139.000 156.600 139.700 156.900 ;
        RECT 140.200 156.600 141.000 157.000 ;
        RECT 131.800 156.200 136.100 156.500 ;
        RECT 136.600 156.500 139.700 156.600 ;
        RECT 136.600 156.300 139.300 156.500 ;
        RECT 136.600 156.200 137.000 156.300 ;
        RECT 125.300 153.400 125.700 155.600 ;
        RECT 126.100 155.300 126.400 156.200 ;
        RECT 126.000 155.000 126.400 155.300 ;
        RECT 129.400 155.000 141.100 155.300 ;
        RECT 126.000 154.000 126.300 155.000 ;
        RECT 129.400 154.700 129.800 155.000 ;
        RECT 138.200 154.800 138.600 155.000 ;
        RECT 140.700 154.900 141.100 155.000 ;
        RECT 126.600 154.300 128.500 154.700 ;
        RECT 126.000 153.700 126.600 154.000 ;
        RECT 120.600 152.800 121.500 153.100 ;
        RECT 123.000 152.800 123.900 153.100 ;
        RECT 125.300 153.000 125.800 153.400 ;
        RECT 118.200 151.100 118.600 152.200 ;
        RECT 121.100 152.200 121.500 152.800 ;
        RECT 123.500 152.200 123.900 152.800 ;
        RECT 121.100 151.800 121.800 152.200 ;
        RECT 123.500 151.800 124.200 152.200 ;
        RECT 121.100 151.100 121.500 151.800 ;
        RECT 123.500 151.100 123.900 151.800 ;
        RECT 125.400 151.100 125.800 153.000 ;
        RECT 126.200 151.100 126.600 153.700 ;
        RECT 128.100 153.700 128.500 154.300 ;
        RECT 128.100 153.400 129.000 153.700 ;
        RECT 128.600 153.100 129.000 153.400 ;
        RECT 131.000 153.200 131.400 154.600 ;
        RECT 132.600 154.300 134.200 154.700 ;
        RECT 136.100 154.300 137.100 154.700 ;
        RECT 141.400 154.500 141.800 157.300 ;
        RECT 143.000 156.000 143.400 159.900 ;
        RECT 144.600 157.600 145.000 159.900 ;
        RECT 132.400 153.900 132.800 154.000 ;
        RECT 132.400 153.600 134.600 153.900 ;
        RECT 134.200 153.500 134.600 153.600 ;
        RECT 135.000 153.400 135.400 154.200 ;
        RECT 128.600 152.700 129.800 153.100 ;
        RECT 131.000 152.800 131.500 153.200 ;
        RECT 133.000 152.800 133.800 153.200 ;
        RECT 134.200 153.100 134.600 153.200 ;
        RECT 136.100 153.100 136.500 154.300 ;
        RECT 137.400 154.100 141.800 154.500 ;
        RECT 139.100 153.400 140.600 153.800 ;
        RECT 139.100 153.100 139.500 153.400 ;
        RECT 134.200 152.800 136.500 153.100 ;
        RECT 129.400 151.100 129.800 152.700 ;
        RECT 138.200 152.700 139.500 153.100 ;
        RECT 130.200 151.100 130.600 152.500 ;
        RECT 131.000 151.100 131.400 152.500 ;
        RECT 131.800 151.100 132.200 152.500 ;
        RECT 132.600 151.100 133.000 152.500 ;
        RECT 134.200 151.100 134.600 152.500 ;
        RECT 135.800 151.100 136.200 152.500 ;
        RECT 136.600 151.100 137.000 152.500 ;
        RECT 137.400 151.100 137.800 152.500 ;
        RECT 138.200 151.100 138.600 152.700 ;
        RECT 141.400 151.100 141.800 154.100 ;
        RECT 142.900 155.600 143.400 156.000 ;
        RECT 143.700 157.300 145.000 157.600 ;
        RECT 143.700 156.500 144.000 157.300 ;
        RECT 146.200 157.200 146.600 159.900 ;
        RECT 147.800 158.500 148.200 159.900 ;
        RECT 148.600 158.500 149.000 159.900 ;
        RECT 149.400 158.500 149.800 159.900 ;
        RECT 146.900 157.200 149.000 157.600 ;
        RECT 145.300 156.800 146.600 157.200 ;
        RECT 150.200 156.800 150.600 159.900 ;
        RECT 151.800 157.500 152.200 159.900 ;
        RECT 153.400 157.500 153.800 159.900 ;
        RECT 154.200 158.500 154.600 159.900 ;
        RECT 155.000 158.500 155.400 159.900 ;
        RECT 156.600 157.600 157.000 159.900 ;
        RECT 158.200 158.200 158.600 159.900 ;
        RECT 162.200 158.200 162.600 159.900 ;
        RECT 158.200 157.900 158.700 158.200 ;
        RECT 158.400 157.600 158.700 157.900 ;
        RECT 162.100 157.900 162.600 158.200 ;
        RECT 162.100 157.600 162.400 157.900 ;
        RECT 163.800 157.600 164.200 159.900 ;
        RECT 165.400 158.500 165.800 159.900 ;
        RECT 166.200 158.500 166.600 159.900 ;
        RECT 156.000 157.200 158.100 157.600 ;
        RECT 158.400 157.300 159.400 157.600 ;
        RECT 151.800 156.800 153.100 157.200 ;
        RECT 153.400 156.900 156.300 157.200 ;
        RECT 157.800 157.000 158.100 157.200 ;
        RECT 147.800 156.500 148.200 156.600 ;
        RECT 143.700 156.200 148.200 156.500 ;
        RECT 149.400 156.500 149.800 156.600 ;
        RECT 153.400 156.500 153.700 156.900 ;
        RECT 156.600 156.600 157.300 156.900 ;
        RECT 157.800 156.600 158.600 157.000 ;
        RECT 149.400 156.200 153.700 156.500 ;
        RECT 154.200 156.500 157.300 156.600 ;
        RECT 154.200 156.300 156.900 156.500 ;
        RECT 154.200 156.200 154.600 156.300 ;
        RECT 142.900 153.400 143.300 155.600 ;
        RECT 143.700 155.300 144.000 156.200 ;
        RECT 158.200 155.800 158.600 156.200 ;
        RECT 158.200 155.300 158.500 155.800 ;
        RECT 143.600 155.000 144.000 155.300 ;
        RECT 147.000 155.000 158.700 155.300 ;
        RECT 143.600 154.000 143.900 155.000 ;
        RECT 147.000 154.700 147.400 155.000 ;
        RECT 155.800 154.800 156.200 155.000 ;
        RECT 158.200 154.900 158.700 155.000 ;
        RECT 158.200 154.800 158.500 154.900 ;
        RECT 144.200 154.300 146.100 154.700 ;
        RECT 143.600 153.700 144.200 154.000 ;
        RECT 142.900 153.000 143.400 153.400 ;
        RECT 143.000 151.100 143.400 153.000 ;
        RECT 143.800 151.100 144.200 153.700 ;
        RECT 145.700 153.700 146.100 154.300 ;
        RECT 145.700 153.400 146.600 153.700 ;
        RECT 146.200 153.100 146.600 153.400 ;
        RECT 148.600 153.200 149.000 154.600 ;
        RECT 150.200 154.300 151.800 154.700 ;
        RECT 153.700 154.300 154.700 154.700 ;
        RECT 159.000 154.500 159.400 157.300 ;
        RECT 150.000 153.900 150.400 154.000 ;
        RECT 150.000 153.600 152.200 153.900 ;
        RECT 151.800 153.500 152.200 153.600 ;
        RECT 152.600 153.400 153.000 154.200 ;
        RECT 146.200 152.700 147.400 153.100 ;
        RECT 148.600 152.800 149.100 153.200 ;
        RECT 150.600 152.800 151.400 153.200 ;
        RECT 151.800 153.100 152.200 153.200 ;
        RECT 153.700 153.100 154.100 154.300 ;
        RECT 155.000 154.100 159.400 154.500 ;
        RECT 156.700 153.400 158.200 153.800 ;
        RECT 156.700 153.100 157.100 153.400 ;
        RECT 151.800 152.800 154.100 153.100 ;
        RECT 147.000 151.100 147.400 152.700 ;
        RECT 155.800 152.700 157.100 153.100 ;
        RECT 147.800 151.100 148.200 152.500 ;
        RECT 148.600 151.100 149.000 152.500 ;
        RECT 149.400 151.100 149.800 152.500 ;
        RECT 150.200 151.100 150.600 152.500 ;
        RECT 151.800 151.100 152.200 152.500 ;
        RECT 153.400 151.100 153.800 152.500 ;
        RECT 154.200 151.100 154.600 152.500 ;
        RECT 155.000 151.100 155.400 152.500 ;
        RECT 155.800 151.100 156.200 152.700 ;
        RECT 159.000 151.100 159.400 154.100 ;
        RECT 161.400 157.300 162.400 157.600 ;
        RECT 161.400 154.500 161.800 157.300 ;
        RECT 162.700 157.200 164.800 157.600 ;
        RECT 167.000 157.500 167.400 159.900 ;
        RECT 168.600 157.500 169.000 159.900 ;
        RECT 162.700 157.000 163.000 157.200 ;
        RECT 162.200 156.600 163.000 157.000 ;
        RECT 164.500 156.900 167.400 157.200 ;
        RECT 163.500 156.600 164.200 156.900 ;
        RECT 163.500 156.500 166.600 156.600 ;
        RECT 163.900 156.300 166.600 156.500 ;
        RECT 166.200 156.200 166.600 156.300 ;
        RECT 167.100 156.500 167.400 156.900 ;
        RECT 167.700 156.800 169.000 157.200 ;
        RECT 170.200 156.800 170.600 159.900 ;
        RECT 171.000 158.500 171.400 159.900 ;
        RECT 171.800 158.500 172.200 159.900 ;
        RECT 172.600 158.500 173.000 159.900 ;
        RECT 171.800 157.200 173.900 157.600 ;
        RECT 174.200 157.200 174.600 159.900 ;
        RECT 175.800 157.600 176.200 159.900 ;
        RECT 175.800 157.300 177.100 157.600 ;
        RECT 174.200 156.800 175.500 157.200 ;
        RECT 171.000 156.500 171.400 156.600 ;
        RECT 167.100 156.200 171.400 156.500 ;
        RECT 172.600 156.500 173.000 156.600 ;
        RECT 176.800 156.500 177.100 157.300 ;
        RECT 172.600 156.200 177.100 156.500 ;
        RECT 176.800 155.300 177.100 156.200 ;
        RECT 177.400 156.000 177.800 159.900 ;
        RECT 179.300 159.200 179.700 159.900 ;
        RECT 179.300 158.800 180.200 159.200 ;
        RECT 179.300 156.300 179.700 158.800 ;
        RECT 181.700 156.300 182.100 159.900 ;
        RECT 177.400 155.600 177.900 156.000 ;
        RECT 179.300 155.900 180.200 156.300 ;
        RECT 181.700 155.900 182.600 156.300 ;
        RECT 185.100 156.200 185.500 159.900 ;
        RECT 162.100 155.000 173.800 155.300 ;
        RECT 176.800 155.000 177.200 155.300 ;
        RECT 162.100 154.900 162.500 155.000 ;
        RECT 163.000 154.800 163.400 155.000 ;
        RECT 164.600 154.800 165.000 155.000 ;
        RECT 173.400 154.700 173.800 155.000 ;
        RECT 161.400 154.100 165.800 154.500 ;
        RECT 166.100 154.300 167.100 154.700 ;
        RECT 169.000 154.300 170.600 154.700 ;
        RECT 161.400 151.100 161.800 154.100 ;
        RECT 162.600 153.400 164.100 153.800 ;
        RECT 163.700 153.100 164.100 153.400 ;
        RECT 166.700 153.100 167.100 154.300 ;
        RECT 167.800 153.400 168.200 154.200 ;
        RECT 170.400 153.900 170.800 154.000 ;
        RECT 168.600 153.600 170.800 153.900 ;
        RECT 168.600 153.500 169.000 153.600 ;
        RECT 171.800 153.200 172.200 154.600 ;
        RECT 174.700 154.300 176.600 154.700 ;
        RECT 174.700 153.700 175.100 154.300 ;
        RECT 176.900 154.000 177.200 155.000 ;
        RECT 168.600 153.100 169.000 153.200 ;
        RECT 163.700 152.700 165.000 153.100 ;
        RECT 166.700 152.800 169.000 153.100 ;
        RECT 169.400 152.800 170.200 153.200 ;
        RECT 171.700 152.800 172.200 153.200 ;
        RECT 174.200 153.400 175.100 153.700 ;
        RECT 176.600 153.700 177.200 154.000 ;
        RECT 174.200 153.100 174.600 153.400 ;
        RECT 164.600 151.100 165.000 152.700 ;
        RECT 173.400 152.700 174.600 153.100 ;
        RECT 165.400 151.100 165.800 152.500 ;
        RECT 166.200 151.100 166.600 152.500 ;
        RECT 167.000 151.100 167.400 152.500 ;
        RECT 168.600 151.100 169.000 152.500 ;
        RECT 170.200 151.100 170.600 152.500 ;
        RECT 171.000 151.100 171.400 152.500 ;
        RECT 171.800 151.100 172.200 152.500 ;
        RECT 172.600 151.100 173.000 152.500 ;
        RECT 173.400 151.100 173.800 152.700 ;
        RECT 176.600 151.100 177.000 153.700 ;
        RECT 177.500 153.400 177.900 155.600 ;
        RECT 179.000 154.800 179.400 155.600 ;
        RECT 179.800 155.100 180.100 155.900 ;
        RECT 181.400 155.100 181.800 155.600 ;
        RECT 179.800 154.800 181.800 155.100 ;
        RECT 177.400 153.000 177.900 153.400 ;
        RECT 179.800 154.200 180.100 154.800 ;
        RECT 182.200 154.200 182.500 155.900 ;
        RECT 184.600 155.800 185.600 156.200 ;
        RECT 184.600 154.400 185.000 155.200 ;
        RECT 185.300 154.200 185.600 155.800 ;
        RECT 179.800 153.800 180.200 154.200 ;
        RECT 182.200 153.800 182.600 154.200 ;
        RECT 183.800 154.100 184.200 154.200 ;
        RECT 183.800 153.800 184.600 154.100 ;
        RECT 185.300 153.800 186.600 154.200 ;
        RECT 177.400 151.100 177.800 153.000 ;
        RECT 179.800 152.100 180.100 153.800 ;
        RECT 180.600 152.400 181.000 153.200 ;
        RECT 182.200 152.200 182.500 153.800 ;
        RECT 184.200 153.600 184.600 153.800 ;
        RECT 183.000 152.400 183.400 153.200 ;
        RECT 183.900 153.100 185.700 153.300 ;
        RECT 186.200 153.100 186.500 153.800 ;
        RECT 183.800 153.000 185.800 153.100 ;
        RECT 179.800 151.100 180.200 152.100 ;
        RECT 182.200 151.100 182.600 152.200 ;
        RECT 183.800 151.100 184.200 153.000 ;
        RECT 185.400 151.100 185.800 153.000 ;
        RECT 186.200 151.100 186.600 153.100 ;
        RECT 187.800 151.100 188.200 159.900 ;
        RECT 189.900 156.200 190.300 159.900 ;
        RECT 189.900 155.900 190.400 156.200 ;
        RECT 190.100 155.200 190.400 155.900 ;
        RECT 191.800 155.900 192.200 159.900 ;
        RECT 193.400 157.900 193.800 159.900 ;
        RECT 191.800 155.200 192.100 155.900 ;
        RECT 193.400 155.800 193.700 157.900 ;
        RECT 192.500 155.500 193.700 155.800 ;
        RECT 195.000 155.700 195.400 159.900 ;
        RECT 197.200 158.200 197.600 159.900 ;
        RECT 196.600 157.900 197.600 158.200 ;
        RECT 199.400 157.900 199.800 159.900 ;
        RECT 201.500 157.900 202.100 159.900 ;
        RECT 196.600 157.500 197.000 157.900 ;
        RECT 199.400 157.600 199.700 157.900 ;
        RECT 198.300 157.300 200.100 157.600 ;
        RECT 201.400 157.500 201.800 157.900 ;
        RECT 198.300 157.200 198.700 157.300 ;
        RECT 199.700 157.200 200.100 157.300 ;
        RECT 196.600 156.500 197.000 156.600 ;
        RECT 198.900 156.500 199.300 156.600 ;
        RECT 196.600 156.200 199.300 156.500 ;
        RECT 199.600 156.500 200.700 156.800 ;
        RECT 199.600 155.900 199.900 156.500 ;
        RECT 200.300 156.400 200.700 156.500 ;
        RECT 201.500 156.600 202.200 157.000 ;
        RECT 201.500 156.100 201.800 156.600 ;
        RECT 197.500 155.700 199.900 155.900 ;
        RECT 195.000 155.600 199.900 155.700 ;
        RECT 200.600 155.800 201.800 156.100 ;
        RECT 195.000 155.500 197.900 155.600 ;
        RECT 189.400 154.400 189.800 155.200 ;
        RECT 190.100 154.800 190.600 155.200 ;
        RECT 191.800 154.800 192.200 155.200 ;
        RECT 190.100 154.200 190.400 154.800 ;
        RECT 188.600 154.100 189.000 154.200 ;
        RECT 188.600 153.800 189.400 154.100 ;
        RECT 190.100 153.800 191.400 154.200 ;
        RECT 189.000 153.600 189.400 153.800 ;
        RECT 188.700 153.100 190.500 153.300 ;
        RECT 191.000 153.100 191.300 153.800 ;
        RECT 191.800 153.100 192.100 154.800 ;
        RECT 192.500 153.800 192.800 155.500 ;
        RECT 195.000 155.400 197.800 155.500 ;
        RECT 198.200 155.100 198.600 155.200 ;
        RECT 196.100 154.800 198.600 155.100 ;
        RECT 196.100 154.700 196.500 154.800 ;
        RECT 194.200 153.800 194.600 154.600 ;
        RECT 196.900 154.200 197.300 154.300 ;
        RECT 200.600 154.200 200.900 155.800 ;
        RECT 203.800 155.600 204.200 159.900 ;
        RECT 202.100 155.300 204.200 155.600 ;
        RECT 202.100 155.200 202.500 155.300 ;
        RECT 202.900 154.900 203.300 155.000 ;
        RECT 201.400 154.600 203.300 154.900 ;
        RECT 201.400 154.500 201.800 154.600 ;
        RECT 195.400 153.900 200.900 154.200 ;
        RECT 195.400 153.800 196.200 153.900 ;
        RECT 192.400 153.700 192.800 153.800 ;
        RECT 192.400 153.500 193.900 153.700 ;
        RECT 192.400 153.400 194.500 153.500 ;
        RECT 193.600 153.200 194.500 153.400 ;
        RECT 194.200 153.100 194.500 153.200 ;
        RECT 188.600 153.000 190.600 153.100 ;
        RECT 188.600 151.100 189.000 153.000 ;
        RECT 190.200 151.100 190.600 153.000 ;
        RECT 191.000 151.100 191.400 153.100 ;
        RECT 191.800 152.600 192.500 153.100 ;
        RECT 192.100 152.200 192.500 152.600 ;
        RECT 191.800 151.800 192.500 152.200 ;
        RECT 192.100 151.100 192.500 151.800 ;
        RECT 194.200 151.100 194.600 153.100 ;
        RECT 195.000 151.100 195.400 153.500 ;
        RECT 197.500 152.800 197.800 153.900 ;
        RECT 200.300 153.800 200.700 153.900 ;
        RECT 203.800 153.600 204.200 155.300 ;
        RECT 202.300 153.300 204.200 153.600 ;
        RECT 202.300 153.200 202.700 153.300 ;
        RECT 196.600 152.100 197.000 152.500 ;
        RECT 197.400 152.400 197.800 152.800 ;
        RECT 198.300 152.700 198.700 152.800 ;
        RECT 198.300 152.400 199.700 152.700 ;
        RECT 199.400 152.100 199.700 152.400 ;
        RECT 201.400 152.100 201.800 152.500 ;
        RECT 196.600 151.800 197.600 152.100 ;
        RECT 197.200 151.100 197.600 151.800 ;
        RECT 199.400 151.100 199.800 152.100 ;
        RECT 201.400 151.800 202.100 152.100 ;
        RECT 201.500 151.100 202.100 151.800 ;
        RECT 203.800 151.100 204.200 153.300 ;
        RECT 0.600 147.500 1.000 149.900 ;
        RECT 2.800 149.200 3.200 149.900 ;
        RECT 2.200 148.900 3.200 149.200 ;
        RECT 5.000 148.900 5.400 149.900 ;
        RECT 7.100 149.200 7.700 149.900 ;
        RECT 7.000 148.900 7.700 149.200 ;
        RECT 2.200 148.500 2.600 148.900 ;
        RECT 5.000 148.600 5.300 148.900 ;
        RECT 3.000 148.200 3.400 148.600 ;
        RECT 3.900 148.300 5.300 148.600 ;
        RECT 7.000 148.500 7.400 148.900 ;
        RECT 3.900 148.200 4.300 148.300 ;
        RECT 3.100 147.200 3.400 148.200 ;
        RECT 7.900 147.700 8.300 147.800 ;
        RECT 9.400 147.700 9.800 149.900 ;
        RECT 10.200 148.000 10.600 149.900 ;
        RECT 11.800 148.000 12.200 149.900 ;
        RECT 10.200 147.900 12.200 148.000 ;
        RECT 12.600 147.900 13.000 149.900 ;
        RECT 15.000 147.900 15.400 149.900 ;
        RECT 15.700 148.200 16.100 148.600 ;
        RECT 17.900 148.200 18.300 149.900 ;
        RECT 10.300 147.700 12.100 147.900 ;
        RECT 7.900 147.400 9.800 147.700 ;
        RECT 1.000 147.100 1.800 147.200 ;
        RECT 3.000 147.100 3.400 147.200 ;
        RECT 5.900 147.100 6.300 147.200 ;
        RECT 1.000 146.800 6.500 147.100 ;
        RECT 2.500 146.700 2.900 146.800 ;
        RECT 1.700 146.200 2.100 146.300 ;
        RECT 6.200 146.200 6.500 146.800 ;
        RECT 7.000 146.400 7.400 146.500 ;
        RECT 1.700 145.900 4.200 146.200 ;
        RECT 3.800 145.800 4.200 145.900 ;
        RECT 6.200 145.800 6.600 146.200 ;
        RECT 7.000 146.100 8.900 146.400 ;
        RECT 8.500 146.000 8.900 146.100 ;
        RECT 0.600 145.500 3.400 145.600 ;
        RECT 0.600 145.400 3.500 145.500 ;
        RECT 0.600 145.300 5.500 145.400 ;
        RECT 0.600 141.100 1.000 145.300 ;
        RECT 3.100 145.100 5.500 145.300 ;
        RECT 2.200 144.500 4.900 144.800 ;
        RECT 2.200 144.400 2.600 144.500 ;
        RECT 4.500 144.400 4.900 144.500 ;
        RECT 5.200 144.500 5.500 145.100 ;
        RECT 6.200 145.200 6.500 145.800 ;
        RECT 7.700 145.700 8.100 145.800 ;
        RECT 9.400 145.700 9.800 147.400 ;
        RECT 10.600 147.200 11.000 147.400 ;
        RECT 12.600 147.200 12.900 147.900 ;
        RECT 10.200 146.900 11.000 147.200 ;
        RECT 10.200 146.800 10.600 146.900 ;
        RECT 11.700 146.800 13.000 147.200 ;
        RECT 13.400 147.100 13.800 147.200 ;
        RECT 14.200 147.100 14.600 147.200 ;
        RECT 13.400 146.800 14.600 147.100 ;
        RECT 11.000 145.800 11.400 146.600 ;
        RECT 7.700 145.400 9.800 145.700 ;
        RECT 6.200 144.900 7.400 145.200 ;
        RECT 5.900 144.500 6.300 144.600 ;
        RECT 5.200 144.200 6.300 144.500 ;
        RECT 7.100 144.400 7.400 144.900 ;
        RECT 7.100 144.000 7.800 144.400 ;
        RECT 3.900 143.700 4.300 143.800 ;
        RECT 5.300 143.700 5.700 143.800 ;
        RECT 2.200 143.100 2.600 143.500 ;
        RECT 3.900 143.400 5.700 143.700 ;
        RECT 5.000 143.100 5.300 143.400 ;
        RECT 7.000 143.100 7.400 143.500 ;
        RECT 2.200 142.800 3.200 143.100 ;
        RECT 2.800 141.100 3.200 142.800 ;
        RECT 5.000 141.100 5.400 143.100 ;
        RECT 7.100 141.100 7.700 143.100 ;
        RECT 9.400 141.100 9.800 145.400 ;
        RECT 11.700 145.100 12.000 146.800 ;
        RECT 14.200 146.400 14.600 146.800 ;
        RECT 13.400 146.100 13.800 146.200 ;
        RECT 15.000 146.100 15.300 147.900 ;
        RECT 15.800 147.800 16.200 148.200 ;
        RECT 17.400 147.900 18.300 148.200 ;
        RECT 19.000 147.900 19.400 149.900 ;
        RECT 19.800 148.000 20.200 149.900 ;
        RECT 21.400 148.000 21.800 149.900 ;
        RECT 19.800 147.900 21.800 148.000 ;
        RECT 16.600 146.800 17.000 147.600 ;
        RECT 17.400 147.100 17.800 147.900 ;
        RECT 19.100 147.200 19.400 147.900 ;
        RECT 19.900 147.700 21.700 147.900 ;
        RECT 22.200 147.500 22.600 149.900 ;
        RECT 24.400 149.200 24.800 149.900 ;
        RECT 23.800 148.900 24.800 149.200 ;
        RECT 26.600 148.900 27.000 149.900 ;
        RECT 28.700 149.200 29.300 149.900 ;
        RECT 28.600 148.900 29.300 149.200 ;
        RECT 23.800 148.500 24.200 148.900 ;
        RECT 26.600 148.600 26.900 148.900 ;
        RECT 24.600 148.200 25.000 148.600 ;
        RECT 25.500 148.300 26.900 148.600 ;
        RECT 28.600 148.500 29.000 148.900 ;
        RECT 25.500 148.200 25.900 148.300 ;
        RECT 21.000 147.200 21.400 147.400 ;
        RECT 18.200 147.100 18.600 147.200 ;
        RECT 17.400 146.800 18.600 147.100 ;
        RECT 19.000 146.800 20.300 147.200 ;
        RECT 21.000 146.900 21.800 147.200 ;
        RECT 21.400 146.800 21.800 146.900 ;
        RECT 22.600 147.100 23.400 147.200 ;
        RECT 24.700 147.100 25.000 148.200 ;
        RECT 29.500 147.700 29.900 147.800 ;
        RECT 31.000 147.700 31.400 149.900 ;
        RECT 29.500 147.400 31.400 147.700 ;
        RECT 31.800 147.500 32.200 149.900 ;
        RECT 34.000 149.200 34.400 149.900 ;
        RECT 33.400 148.900 34.400 149.200 ;
        RECT 36.200 148.900 36.600 149.900 ;
        RECT 38.300 149.200 38.900 149.900 ;
        RECT 38.200 148.900 38.900 149.200 ;
        RECT 33.400 148.500 33.800 148.900 ;
        RECT 36.200 148.600 36.500 148.900 ;
        RECT 34.200 148.200 34.600 148.600 ;
        RECT 35.100 148.300 36.500 148.600 ;
        RECT 38.200 148.500 38.600 148.900 ;
        RECT 35.100 148.200 35.500 148.300 ;
        RECT 27.500 147.100 27.900 147.200 ;
        RECT 22.600 146.800 28.100 147.100 ;
        RECT 15.800 146.100 16.200 146.200 ;
        RECT 13.400 145.800 14.200 146.100 ;
        RECT 15.000 145.800 16.200 146.100 ;
        RECT 13.800 145.600 14.200 145.800 ;
        RECT 12.600 145.100 13.000 145.200 ;
        RECT 15.800 145.100 16.100 145.800 ;
        RECT 11.500 144.800 12.000 145.100 ;
        RECT 12.300 144.800 13.000 145.100 ;
        RECT 13.400 144.800 15.400 145.100 ;
        RECT 11.500 141.100 11.900 144.800 ;
        RECT 12.300 144.200 12.600 144.800 ;
        RECT 12.200 143.800 12.600 144.200 ;
        RECT 13.400 141.100 13.800 144.800 ;
        RECT 15.000 141.100 15.400 144.800 ;
        RECT 15.800 141.100 16.200 145.100 ;
        RECT 17.400 141.100 17.800 146.800 ;
        RECT 18.200 144.400 18.600 145.200 ;
        RECT 19.000 145.100 19.400 145.200 ;
        RECT 20.000 145.100 20.300 146.800 ;
        RECT 24.100 146.700 24.500 146.800 ;
        RECT 20.600 145.800 21.000 146.600 ;
        RECT 23.300 146.200 23.700 146.300 ;
        RECT 24.600 146.200 25.000 146.300 ;
        RECT 23.300 145.900 25.800 146.200 ;
        RECT 25.400 145.800 25.800 145.900 ;
        RECT 22.200 145.500 25.000 145.600 ;
        RECT 22.200 145.400 25.100 145.500 ;
        RECT 22.200 145.300 27.100 145.400 ;
        RECT 19.000 144.800 19.700 145.100 ;
        RECT 20.000 144.800 20.500 145.100 ;
        RECT 19.400 144.200 19.700 144.800 ;
        RECT 19.400 143.800 19.800 144.200 ;
        RECT 20.100 141.100 20.500 144.800 ;
        RECT 22.200 141.100 22.600 145.300 ;
        RECT 24.700 145.100 27.100 145.300 ;
        RECT 23.800 144.500 26.500 144.800 ;
        RECT 23.800 144.400 24.200 144.500 ;
        RECT 26.100 144.400 26.500 144.500 ;
        RECT 26.800 144.500 27.100 145.100 ;
        RECT 27.800 145.200 28.100 146.800 ;
        RECT 28.600 146.400 29.000 146.500 ;
        RECT 28.600 146.100 30.500 146.400 ;
        RECT 30.100 146.000 30.500 146.100 ;
        RECT 29.300 145.700 29.700 145.800 ;
        RECT 31.000 145.700 31.400 147.400 ;
        RECT 32.200 147.100 33.000 147.200 ;
        RECT 34.300 147.100 34.600 148.200 ;
        RECT 39.100 147.700 39.500 147.800 ;
        RECT 40.600 147.700 41.000 149.900 ;
        RECT 39.100 147.400 41.000 147.700 ;
        RECT 41.400 147.500 41.800 149.900 ;
        RECT 43.600 149.200 44.000 149.900 ;
        RECT 43.000 148.900 44.000 149.200 ;
        RECT 45.800 148.900 46.200 149.900 ;
        RECT 47.900 149.200 48.500 149.900 ;
        RECT 47.800 148.900 48.500 149.200 ;
        RECT 43.000 148.500 43.400 148.900 ;
        RECT 45.800 148.600 46.100 148.900 ;
        RECT 43.800 148.200 44.200 148.600 ;
        RECT 44.700 148.300 46.100 148.600 ;
        RECT 47.800 148.500 48.200 148.900 ;
        RECT 44.700 148.200 45.100 148.300 ;
        RECT 35.800 147.100 36.200 147.200 ;
        RECT 37.100 147.100 37.500 147.200 ;
        RECT 32.200 146.800 37.700 147.100 ;
        RECT 39.800 146.800 40.200 147.400 ;
        RECT 33.700 146.700 34.100 146.800 ;
        RECT 32.900 146.200 33.300 146.300 ;
        RECT 32.900 146.100 35.400 146.200 ;
        RECT 36.600 146.100 37.000 146.200 ;
        RECT 32.900 145.900 37.000 146.100 ;
        RECT 35.000 145.800 37.000 145.900 ;
        RECT 29.300 145.400 31.400 145.700 ;
        RECT 27.800 144.900 29.000 145.200 ;
        RECT 27.500 144.500 27.900 144.600 ;
        RECT 26.800 144.200 27.900 144.500 ;
        RECT 28.700 144.400 29.000 144.900 ;
        RECT 28.700 144.000 29.400 144.400 ;
        RECT 25.500 143.700 25.900 143.800 ;
        RECT 26.900 143.700 27.300 143.800 ;
        RECT 23.800 143.100 24.200 143.500 ;
        RECT 25.500 143.400 27.300 143.700 ;
        RECT 26.600 143.100 26.900 143.400 ;
        RECT 28.600 143.100 29.000 143.500 ;
        RECT 23.800 142.800 24.800 143.100 ;
        RECT 24.400 141.100 24.800 142.800 ;
        RECT 26.600 141.100 27.000 143.100 ;
        RECT 28.700 141.100 29.300 143.100 ;
        RECT 31.000 141.100 31.400 145.400 ;
        RECT 31.800 145.500 34.600 145.600 ;
        RECT 31.800 145.400 34.700 145.500 ;
        RECT 31.800 145.300 36.700 145.400 ;
        RECT 31.800 141.100 32.200 145.300 ;
        RECT 34.300 145.100 36.700 145.300 ;
        RECT 33.400 144.500 36.100 144.800 ;
        RECT 33.400 144.400 33.800 144.500 ;
        RECT 35.700 144.400 36.100 144.500 ;
        RECT 36.400 144.500 36.700 145.100 ;
        RECT 37.400 145.200 37.700 146.800 ;
        RECT 38.200 146.400 38.600 146.500 ;
        RECT 38.200 146.100 40.100 146.400 ;
        RECT 39.700 146.000 40.100 146.100 ;
        RECT 38.900 145.700 39.300 145.800 ;
        RECT 40.600 145.700 41.000 147.400 ;
        RECT 41.800 147.100 42.600 147.200 ;
        RECT 43.900 147.100 44.200 148.200 ;
        RECT 48.700 147.700 49.100 147.800 ;
        RECT 50.200 147.700 50.600 149.900 ;
        RECT 48.700 147.400 50.600 147.700 ;
        RECT 44.600 147.100 45.000 147.200 ;
        RECT 46.700 147.100 47.100 147.200 ;
        RECT 41.800 146.800 47.300 147.100 ;
        RECT 43.300 146.700 43.700 146.800 ;
        RECT 42.500 146.200 42.900 146.300 ;
        RECT 42.500 146.100 45.000 146.200 ;
        RECT 46.200 146.100 46.600 146.200 ;
        RECT 42.500 145.900 46.600 146.100 ;
        RECT 44.600 145.800 46.600 145.900 ;
        RECT 38.900 145.400 41.000 145.700 ;
        RECT 37.400 144.900 38.600 145.200 ;
        RECT 37.100 144.500 37.500 144.600 ;
        RECT 36.400 144.200 37.500 144.500 ;
        RECT 38.300 144.400 38.600 144.900 ;
        RECT 38.300 144.000 39.000 144.400 ;
        RECT 35.100 143.700 35.500 143.800 ;
        RECT 36.500 143.700 36.900 143.800 ;
        RECT 33.400 143.100 33.800 143.500 ;
        RECT 35.100 143.400 36.900 143.700 ;
        RECT 36.200 143.100 36.500 143.400 ;
        RECT 38.200 143.100 38.600 143.500 ;
        RECT 33.400 142.800 34.400 143.100 ;
        RECT 34.000 141.100 34.400 142.800 ;
        RECT 36.200 141.100 36.600 143.100 ;
        RECT 38.300 141.100 38.900 143.100 ;
        RECT 40.600 141.100 41.000 145.400 ;
        RECT 41.400 145.500 44.200 145.600 ;
        RECT 41.400 145.400 44.300 145.500 ;
        RECT 41.400 145.300 46.300 145.400 ;
        RECT 41.400 141.100 41.800 145.300 ;
        RECT 43.900 145.100 46.300 145.300 ;
        RECT 43.000 144.500 45.700 144.800 ;
        RECT 43.000 144.400 43.400 144.500 ;
        RECT 45.300 144.400 45.700 144.500 ;
        RECT 46.000 144.500 46.300 145.100 ;
        RECT 47.000 145.200 47.300 146.800 ;
        RECT 47.800 146.400 48.200 146.500 ;
        RECT 47.800 146.100 49.700 146.400 ;
        RECT 49.300 146.000 49.700 146.100 ;
        RECT 48.500 145.700 48.900 145.800 ;
        RECT 50.200 145.700 50.600 147.400 ;
        RECT 48.500 145.400 50.600 145.700 ;
        RECT 47.000 144.900 48.200 145.200 ;
        RECT 46.700 144.500 47.100 144.600 ;
        RECT 46.000 144.200 47.100 144.500 ;
        RECT 47.900 144.400 48.200 144.900 ;
        RECT 47.900 144.000 48.600 144.400 ;
        RECT 44.700 143.700 45.100 143.800 ;
        RECT 46.100 143.700 46.500 143.800 ;
        RECT 43.000 143.100 43.400 143.500 ;
        RECT 44.700 143.400 46.500 143.700 ;
        RECT 45.800 143.100 46.100 143.400 ;
        RECT 47.800 143.100 48.200 143.500 ;
        RECT 43.000 142.800 44.000 143.100 ;
        RECT 43.600 141.100 44.000 142.800 ;
        RECT 45.800 141.100 46.200 143.100 ;
        RECT 47.900 141.100 48.500 143.100 ;
        RECT 50.200 142.100 50.600 145.400 ;
        RECT 51.800 142.100 52.200 142.200 ;
        RECT 50.200 141.800 52.200 142.100 ;
        RECT 50.200 141.100 50.600 141.800 ;
        RECT 52.600 141.100 53.000 149.900 ;
        RECT 53.400 147.800 53.800 148.600 ;
        RECT 55.500 148.200 55.900 149.900 ;
        RECT 55.000 147.900 55.900 148.200 ;
        RECT 56.600 147.900 57.000 149.900 ;
        RECT 57.400 148.000 57.800 149.900 ;
        RECT 59.000 148.000 59.400 149.900 ;
        RECT 57.400 147.900 59.400 148.000 ;
        RECT 54.200 146.800 54.600 147.600 ;
        RECT 55.000 146.100 55.400 147.900 ;
        RECT 56.700 147.200 57.000 147.900 ;
        RECT 57.500 147.700 59.300 147.900 ;
        RECT 59.800 147.600 60.200 149.900 ;
        RECT 61.400 148.200 61.800 149.900 ;
        RECT 61.400 147.900 61.900 148.200 ;
        RECT 58.600 147.200 59.000 147.400 ;
        RECT 59.800 147.300 61.100 147.600 ;
        RECT 56.600 146.800 57.900 147.200 ;
        RECT 58.600 146.900 59.400 147.200 ;
        RECT 59.000 146.800 59.400 146.900 ;
        RECT 55.000 145.800 56.900 146.100 ;
        RECT 55.000 141.100 55.400 145.800 ;
        RECT 56.600 145.200 56.900 145.800 ;
        RECT 55.800 144.400 56.200 145.200 ;
        RECT 56.600 145.100 57.000 145.200 ;
        RECT 57.600 145.100 57.900 146.800 ;
        RECT 58.200 145.800 58.600 146.600 ;
        RECT 59.900 146.200 60.300 146.600 ;
        RECT 59.800 145.800 60.300 146.200 ;
        RECT 60.800 146.500 61.100 147.300 ;
        RECT 61.600 147.200 61.900 147.900 ;
        RECT 63.000 147.800 63.400 148.600 ;
        RECT 61.400 146.800 61.900 147.200 ;
        RECT 60.800 146.100 61.300 146.500 ;
        RECT 60.800 145.100 61.100 146.100 ;
        RECT 61.600 145.100 61.900 146.800 ;
        RECT 56.600 144.800 57.300 145.100 ;
        RECT 57.600 144.800 58.100 145.100 ;
        RECT 57.000 144.200 57.300 144.800 ;
        RECT 57.000 143.800 57.400 144.200 ;
        RECT 57.700 141.100 58.100 144.800 ;
        RECT 59.800 144.800 61.100 145.100 ;
        RECT 59.800 141.100 60.200 144.800 ;
        RECT 61.400 144.600 61.900 145.100 ;
        RECT 61.400 141.100 61.800 144.600 ;
        RECT 63.800 141.100 64.200 149.900 ;
        RECT 65.400 148.800 65.800 149.900 ;
        RECT 65.400 147.200 65.700 148.800 ;
        RECT 66.200 148.100 66.600 148.600 ;
        RECT 67.000 148.100 67.400 148.200 ;
        RECT 66.200 147.800 67.400 148.100 ;
        RECT 67.800 148.000 68.200 149.900 ;
        RECT 67.700 147.600 68.200 148.000 ;
        RECT 65.400 146.800 65.800 147.200 ;
        RECT 64.600 145.400 65.000 146.200 ;
        RECT 65.400 145.100 65.700 146.800 ;
        RECT 67.700 145.400 68.100 147.600 ;
        RECT 68.600 147.300 69.000 149.900 ;
        RECT 71.800 148.300 72.200 149.900 ;
        RECT 72.600 148.500 73.000 149.900 ;
        RECT 73.400 148.500 73.800 149.900 ;
        RECT 74.200 148.500 74.600 149.900 ;
        RECT 75.000 148.500 75.400 149.900 ;
        RECT 76.600 148.500 77.000 149.900 ;
        RECT 78.200 148.500 78.600 149.900 ;
        RECT 79.000 148.500 79.400 149.900 ;
        RECT 79.800 148.500 80.200 149.900 ;
        RECT 71.000 147.900 72.200 148.300 ;
        RECT 80.600 148.300 81.000 149.900 ;
        RECT 71.000 147.600 71.400 147.900 ;
        RECT 68.400 147.000 69.000 147.300 ;
        RECT 70.500 147.300 71.400 147.600 ;
        RECT 73.400 147.800 73.900 148.200 ;
        RECT 75.400 147.800 76.200 148.200 ;
        RECT 76.600 147.900 78.900 148.200 ;
        RECT 80.600 147.900 81.900 148.300 ;
        RECT 76.600 147.800 77.000 147.900 ;
        RECT 68.400 146.000 68.700 147.000 ;
        RECT 70.500 146.700 70.900 147.300 ;
        RECT 69.000 146.300 70.900 146.700 ;
        RECT 73.400 146.400 73.800 147.800 ;
        RECT 76.600 147.400 77.000 147.500 ;
        RECT 74.800 147.100 77.000 147.400 ;
        RECT 74.800 147.000 75.200 147.100 ;
        RECT 77.400 146.800 77.800 147.600 ;
        RECT 78.500 146.700 78.900 147.900 ;
        RECT 81.500 147.600 81.900 147.900 ;
        RECT 81.500 147.200 83.000 147.600 ;
        RECT 83.800 146.900 84.200 149.900 ;
        RECT 84.600 147.800 85.000 148.600 ;
        RECT 75.000 146.300 76.600 146.700 ;
        RECT 78.500 146.300 79.500 146.700 ;
        RECT 79.800 146.500 84.200 146.900 ;
        RECT 71.800 146.000 72.200 146.300 ;
        RECT 80.600 146.000 81.000 146.200 ;
        RECT 81.400 146.000 81.800 146.200 ;
        RECT 83.100 146.000 83.500 146.100 ;
        RECT 68.400 145.700 68.800 146.000 ;
        RECT 71.800 145.700 83.500 146.000 ;
        RECT 64.900 144.700 65.800 145.100 ;
        RECT 67.700 145.000 68.200 145.400 ;
        RECT 64.900 141.100 65.300 144.700 ;
        RECT 67.800 141.100 68.200 145.000 ;
        RECT 68.500 144.800 68.800 145.700 ;
        RECT 68.500 144.500 73.000 144.800 ;
        RECT 68.500 143.700 68.800 144.500 ;
        RECT 72.600 144.400 73.000 144.500 ;
        RECT 74.200 144.500 78.500 144.800 ;
        RECT 74.200 144.400 74.600 144.500 ;
        RECT 70.100 143.800 71.400 144.200 ;
        RECT 68.500 143.400 69.800 143.700 ;
        RECT 69.400 141.100 69.800 143.400 ;
        RECT 71.000 141.100 71.400 143.800 ;
        RECT 71.700 143.400 73.800 143.800 ;
        RECT 72.600 141.100 73.000 142.500 ;
        RECT 73.400 141.100 73.800 142.500 ;
        RECT 74.200 141.100 74.600 142.500 ;
        RECT 75.000 141.100 75.400 144.200 ;
        RECT 76.600 143.800 77.900 144.200 ;
        RECT 78.200 144.100 78.500 144.500 ;
        RECT 79.000 144.700 79.400 144.800 ;
        RECT 79.000 144.500 81.700 144.700 ;
        RECT 79.000 144.400 82.100 144.500 ;
        RECT 81.400 144.100 82.100 144.400 ;
        RECT 78.200 143.800 81.100 144.100 ;
        RECT 82.600 144.000 83.400 144.400 ;
        RECT 82.600 143.800 82.900 144.000 ;
        RECT 76.600 141.100 77.000 143.500 ;
        RECT 78.200 141.100 78.600 143.500 ;
        RECT 80.800 143.400 82.900 143.800 ;
        RECT 83.800 143.700 84.200 146.500 ;
        RECT 83.200 143.400 84.200 143.700 ;
        RECT 79.000 141.100 79.400 142.500 ;
        RECT 79.800 141.100 80.200 142.500 ;
        RECT 81.400 141.100 81.800 143.400 ;
        RECT 83.200 143.100 83.500 143.400 ;
        RECT 83.000 142.800 83.500 143.100 ;
        RECT 83.000 141.100 83.400 142.800 ;
        RECT 85.400 141.100 85.800 149.900 ;
        RECT 86.200 148.000 86.600 149.900 ;
        RECT 87.800 148.000 88.200 149.900 ;
        RECT 86.200 147.900 88.200 148.000 ;
        RECT 88.600 147.900 89.000 149.900 ;
        RECT 89.700 148.200 90.100 149.900 ;
        RECT 89.700 147.900 90.600 148.200 ;
        RECT 86.300 147.700 88.100 147.900 ;
        RECT 86.600 147.200 87.000 147.400 ;
        RECT 88.600 147.200 88.900 147.900 ;
        RECT 86.200 146.900 87.000 147.200 ;
        RECT 86.200 146.800 86.600 146.900 ;
        RECT 87.700 146.800 89.000 147.200 ;
        RECT 87.000 145.800 87.400 146.600 ;
        RECT 87.700 145.100 88.000 146.800 ;
        RECT 90.200 146.100 90.600 147.900 ;
        RECT 91.800 147.700 92.200 149.900 ;
        RECT 93.900 149.200 94.500 149.900 ;
        RECT 93.900 148.900 94.600 149.200 ;
        RECT 96.200 148.900 96.600 149.900 ;
        RECT 98.400 149.200 98.800 149.900 ;
        RECT 98.400 148.900 99.400 149.200 ;
        RECT 94.200 148.500 94.600 148.900 ;
        RECT 96.300 148.600 96.600 148.900 ;
        RECT 96.300 148.300 97.700 148.600 ;
        RECT 97.300 148.200 97.700 148.300 ;
        RECT 98.200 148.200 98.600 148.600 ;
        RECT 99.000 148.500 99.400 148.900 ;
        RECT 93.300 147.700 93.700 147.800 ;
        RECT 91.000 147.100 91.400 147.600 ;
        RECT 91.800 147.400 93.700 147.700 ;
        RECT 91.800 147.100 92.200 147.400 ;
        RECT 95.300 147.100 95.700 147.200 ;
        RECT 98.200 147.100 98.500 148.200 ;
        RECT 100.600 147.500 101.000 149.900 ;
        RECT 99.800 147.100 100.600 147.200 ;
        RECT 101.400 147.100 101.800 147.200 ;
        RECT 103.600 147.100 104.000 149.900 ;
        RECT 91.000 146.800 92.200 147.100 ;
        RECT 88.600 145.800 90.600 146.100 ;
        RECT 88.600 145.200 88.900 145.800 ;
        RECT 88.600 145.100 89.000 145.200 ;
        RECT 87.500 144.800 88.000 145.100 ;
        RECT 88.300 144.800 89.000 145.100 ;
        RECT 87.500 141.100 87.900 144.800 ;
        RECT 88.300 144.200 88.600 144.800 ;
        RECT 89.400 144.400 89.800 145.200 ;
        RECT 88.200 143.800 88.600 144.200 ;
        RECT 90.200 141.100 90.600 145.800 ;
        RECT 91.800 145.700 92.200 146.800 ;
        RECT 95.100 146.800 101.800 147.100 ;
        RECT 103.100 146.900 104.000 147.100 ;
        RECT 108.000 147.100 108.400 149.900 ;
        RECT 110.200 148.900 110.600 149.900 ;
        RECT 110.200 147.200 110.500 148.900 ;
        RECT 111.000 148.100 111.400 148.600 ;
        RECT 112.100 148.200 112.500 149.900 ;
        RECT 112.100 148.100 113.000 148.200 ;
        RECT 111.000 147.800 113.000 148.100 ;
        RECT 108.000 146.900 108.900 147.100 ;
        RECT 103.100 146.800 103.900 146.900 ;
        RECT 108.100 146.800 108.900 146.900 ;
        RECT 94.200 146.400 94.600 146.500 ;
        RECT 92.700 146.100 94.600 146.400 ;
        RECT 95.100 146.200 95.400 146.800 ;
        RECT 98.700 146.700 99.100 146.800 ;
        RECT 99.500 146.200 99.900 146.300 ;
        RECT 92.700 146.000 93.100 146.100 ;
        RECT 95.000 145.800 95.400 146.200 ;
        RECT 95.800 146.100 96.200 146.200 ;
        RECT 97.400 146.100 99.900 146.200 ;
        RECT 95.800 145.900 99.900 146.100 ;
        RECT 95.800 145.800 97.800 145.900 ;
        RECT 93.500 145.700 93.900 145.800 ;
        RECT 91.800 145.400 93.900 145.700 ;
        RECT 91.800 141.100 92.200 145.400 ;
        RECT 95.100 145.200 95.400 145.800 ;
        RECT 98.200 145.500 101.000 145.600 ;
        RECT 98.100 145.400 101.000 145.500 ;
        RECT 94.200 144.900 95.400 145.200 ;
        RECT 96.100 145.300 101.000 145.400 ;
        RECT 96.100 145.100 98.500 145.300 ;
        RECT 94.200 144.400 94.500 144.900 ;
        RECT 93.800 144.000 94.500 144.400 ;
        RECT 95.300 144.500 95.700 144.600 ;
        RECT 96.100 144.500 96.400 145.100 ;
        RECT 95.300 144.200 96.400 144.500 ;
        RECT 96.700 144.500 99.400 144.800 ;
        RECT 96.700 144.400 97.100 144.500 ;
        RECT 99.000 144.400 99.400 144.500 ;
        RECT 95.900 143.700 96.300 143.800 ;
        RECT 97.300 143.700 97.700 143.800 ;
        RECT 94.200 143.100 94.600 143.500 ;
        RECT 95.900 143.400 97.700 143.700 ;
        RECT 96.300 143.100 96.600 143.400 ;
        RECT 99.000 143.100 99.400 143.500 ;
        RECT 93.900 141.100 94.500 143.100 ;
        RECT 96.200 141.100 96.600 143.100 ;
        RECT 98.400 142.800 99.400 143.100 ;
        RECT 98.400 141.100 98.800 142.800 ;
        RECT 100.600 141.100 101.000 145.300 ;
        RECT 103.100 145.200 103.400 146.800 ;
        RECT 104.200 145.800 105.000 146.200 ;
        RECT 103.000 144.800 103.400 145.200 ;
        RECT 105.400 145.100 105.800 146.200 ;
        RECT 107.000 145.800 107.800 146.200 ;
        RECT 106.200 145.100 106.600 145.600 ;
        RECT 105.400 144.800 106.600 145.100 ;
        RECT 108.600 145.200 108.900 146.800 ;
        RECT 110.200 146.800 110.600 147.200 ;
        RECT 109.400 145.400 109.800 146.200 ;
        RECT 108.600 144.800 109.000 145.200 ;
        RECT 110.200 145.100 110.500 146.800 ;
        RECT 103.100 143.500 103.400 144.800 ;
        RECT 103.800 143.800 104.200 144.600 ;
        RECT 107.000 143.800 107.400 144.200 ;
        RECT 107.800 143.800 108.200 144.600 ;
        RECT 107.000 143.500 107.300 143.800 ;
        RECT 108.600 143.500 108.900 144.800 ;
        RECT 103.100 143.200 104.900 143.500 ;
        RECT 103.100 143.100 103.400 143.200 ;
        RECT 103.000 141.100 103.400 143.100 ;
        RECT 104.600 143.100 104.900 143.200 ;
        RECT 107.000 143.200 108.900 143.500 ;
        RECT 104.600 141.100 105.000 143.100 ;
        RECT 107.000 141.100 107.400 143.200 ;
        RECT 108.600 143.100 108.900 143.200 ;
        RECT 109.700 144.700 110.600 145.100 ;
        RECT 108.600 141.100 109.000 143.100 ;
        RECT 109.700 142.200 110.100 144.700 ;
        RECT 111.800 144.400 112.200 145.200 ;
        RECT 109.400 141.800 110.100 142.200 ;
        RECT 109.700 141.100 110.100 141.800 ;
        RECT 112.600 141.100 113.000 147.800 ;
        RECT 113.400 146.800 113.800 147.600 ;
        RECT 116.000 147.100 116.400 149.900 ;
        RECT 119.200 147.100 119.600 149.900 ;
        RECT 122.400 147.100 122.800 149.900 ;
        RECT 125.600 147.100 126.000 149.900 ;
        RECT 128.800 147.100 129.200 149.900 ;
        RECT 131.000 148.900 131.400 149.900 ;
        RECT 130.200 147.800 130.600 148.600 ;
        RECT 131.100 147.200 131.400 148.900 ;
        RECT 133.400 148.200 133.800 149.900 ;
        RECT 116.000 146.900 116.900 147.100 ;
        RECT 119.200 146.900 120.100 147.100 ;
        RECT 122.400 146.900 123.300 147.100 ;
        RECT 125.600 146.900 126.500 147.100 ;
        RECT 128.800 146.900 129.700 147.100 ;
        RECT 116.100 146.800 116.900 146.900 ;
        RECT 119.300 146.800 120.100 146.900 ;
        RECT 122.500 146.800 123.300 146.900 ;
        RECT 125.700 146.800 126.500 146.900 ;
        RECT 128.900 146.800 129.700 146.900 ;
        RECT 131.000 146.800 131.400 147.200 ;
        RECT 115.000 145.800 115.800 146.200 ;
        RECT 114.200 144.800 114.600 145.600 ;
        RECT 116.600 145.200 116.900 146.800 ;
        RECT 118.200 145.800 119.000 146.200 ;
        RECT 116.600 144.800 117.000 145.200 ;
        RECT 117.400 144.800 117.800 145.600 ;
        RECT 119.800 145.200 120.100 146.800 ;
        RECT 121.400 145.800 122.200 146.200 ;
        RECT 119.800 144.800 120.200 145.200 ;
        RECT 120.600 144.800 121.000 145.600 ;
        RECT 123.000 145.200 123.300 146.800 ;
        RECT 124.600 145.800 125.400 146.200 ;
        RECT 123.000 144.800 123.400 145.200 ;
        RECT 123.800 144.800 124.200 145.600 ;
        RECT 126.200 145.200 126.500 146.800 ;
        RECT 126.200 144.800 126.600 145.200 ;
        RECT 127.000 144.800 127.400 146.200 ;
        RECT 127.800 145.800 128.600 146.200 ;
        RECT 129.400 145.200 129.700 146.800 ;
        RECT 129.400 144.800 129.800 145.200 ;
        RECT 131.100 145.100 131.400 146.800 ;
        RECT 133.300 147.900 133.800 148.200 ;
        RECT 133.300 147.200 133.600 147.900 ;
        RECT 135.000 147.600 135.400 149.900 ;
        RECT 136.600 148.900 137.000 149.900 ;
        RECT 135.800 147.800 136.200 148.600 ;
        RECT 134.100 147.300 135.400 147.600 ;
        RECT 133.300 146.800 133.800 147.200 ;
        RECT 131.800 145.400 132.200 146.200 ;
        RECT 133.300 145.100 133.600 146.800 ;
        RECT 134.100 146.500 134.400 147.300 ;
        RECT 136.700 147.200 137.000 148.900 ;
        RECT 138.200 147.900 138.600 149.900 ;
        RECT 140.400 148.100 141.200 149.900 ;
        RECT 138.200 147.600 139.400 147.900 ;
        RECT 139.000 147.500 139.400 147.600 ;
        RECT 139.700 147.400 140.100 147.800 ;
        RECT 139.700 147.200 140.000 147.400 ;
        RECT 136.600 146.800 137.000 147.200 ;
        RECT 138.200 146.800 139.000 147.200 ;
        RECT 139.600 146.800 140.000 147.200 ;
        RECT 133.900 146.100 134.400 146.500 ;
        RECT 134.100 145.100 134.400 146.100 ;
        RECT 134.900 146.200 135.300 146.600 ;
        RECT 134.900 145.800 135.400 146.200 ;
        RECT 136.700 145.100 137.000 146.800 ;
        RECT 140.400 146.400 140.700 148.100 ;
        RECT 143.000 147.900 143.400 149.900 ;
        RECT 145.100 148.200 145.500 149.900 ;
        RECT 147.500 148.200 147.900 149.900 ;
        RECT 141.000 147.700 141.800 147.800 ;
        RECT 141.000 147.400 142.000 147.700 ;
        RECT 142.300 147.600 143.400 147.900 ;
        RECT 144.600 147.900 145.500 148.200 ;
        RECT 147.000 147.900 147.900 148.200 ;
        RECT 150.200 147.900 150.600 149.900 ;
        RECT 150.900 148.200 151.300 148.600 ;
        RECT 142.300 147.500 142.700 147.600 ;
        RECT 141.700 147.200 142.000 147.400 ;
        RECT 141.000 146.700 141.400 147.100 ;
        RECT 141.700 146.900 143.400 147.200 ;
        RECT 142.600 146.800 143.400 146.900 ;
        RECT 143.800 146.800 144.200 147.600 ;
        RECT 140.200 146.200 140.700 146.400 ;
        RECT 137.400 145.400 137.800 146.200 ;
        RECT 139.800 146.100 140.700 146.200 ;
        RECT 141.100 146.400 141.400 146.700 ;
        RECT 141.100 146.100 142.400 146.400 ;
        RECT 139.800 145.800 140.500 146.100 ;
        RECT 142.000 146.000 142.400 146.100 ;
        RECT 143.000 146.100 143.300 146.800 ;
        RECT 144.600 146.100 145.000 147.900 ;
        RECT 146.200 146.800 146.600 147.600 ;
        RECT 143.000 145.800 145.000 146.100 ;
        RECT 140.200 145.100 140.500 145.800 ;
        RECT 140.900 145.700 141.300 145.800 ;
        RECT 140.900 145.400 142.600 145.700 ;
        RECT 142.300 145.100 142.600 145.400 ;
        RECT 115.800 143.800 116.200 144.600 ;
        RECT 116.600 143.500 116.900 144.800 ;
        RECT 117.400 144.200 117.700 144.800 ;
        RECT 117.400 143.800 117.800 144.200 ;
        RECT 119.000 143.800 119.400 144.600 ;
        RECT 119.800 143.500 120.100 144.800 ;
        RECT 122.200 143.800 122.600 144.600 ;
        RECT 123.000 143.500 123.300 144.800 ;
        RECT 125.400 143.800 125.800 144.600 ;
        RECT 126.200 143.500 126.500 144.800 ;
        RECT 128.600 143.800 129.000 144.600 ;
        RECT 129.400 143.500 129.700 144.800 ;
        RECT 131.000 144.700 131.900 145.100 ;
        RECT 115.100 143.200 116.900 143.500 ;
        RECT 115.100 143.100 115.400 143.200 ;
        RECT 115.000 141.100 115.400 143.100 ;
        RECT 116.600 143.100 116.900 143.200 ;
        RECT 118.300 143.200 120.100 143.500 ;
        RECT 118.300 143.100 118.600 143.200 ;
        RECT 116.600 141.100 117.000 143.100 ;
        RECT 118.200 141.100 118.600 143.100 ;
        RECT 119.800 143.100 120.100 143.200 ;
        RECT 121.500 143.200 123.300 143.500 ;
        RECT 121.500 143.100 121.800 143.200 ;
        RECT 119.800 141.100 120.200 143.100 ;
        RECT 121.400 141.100 121.800 143.100 ;
        RECT 123.000 143.100 123.300 143.200 ;
        RECT 124.700 143.200 126.500 143.500 ;
        RECT 124.700 143.100 125.000 143.200 ;
        RECT 123.000 141.100 123.400 143.100 ;
        RECT 124.600 141.100 125.000 143.100 ;
        RECT 126.200 143.100 126.500 143.200 ;
        RECT 127.900 143.200 129.700 143.500 ;
        RECT 127.900 143.100 128.200 143.200 ;
        RECT 126.200 141.100 126.600 143.100 ;
        RECT 127.800 141.100 128.200 143.100 ;
        RECT 129.400 143.100 129.700 143.200 ;
        RECT 129.400 141.100 129.800 143.100 ;
        RECT 131.500 142.200 131.900 144.700 ;
        RECT 133.300 144.600 133.800 145.100 ;
        RECT 134.100 144.800 135.400 145.100 ;
        RECT 131.000 141.800 131.900 142.200 ;
        RECT 131.500 141.100 131.900 141.800 ;
        RECT 133.400 141.100 133.800 144.600 ;
        RECT 135.000 141.100 135.400 144.800 ;
        RECT 136.600 144.700 137.500 145.100 ;
        RECT 137.100 141.100 137.500 144.700 ;
        RECT 138.200 144.800 139.400 145.100 ;
        RECT 140.200 144.800 141.200 145.100 ;
        RECT 138.200 141.100 138.600 144.800 ;
        RECT 139.000 144.700 139.400 144.800 ;
        RECT 140.400 141.100 141.200 144.800 ;
        RECT 142.300 144.800 143.400 145.100 ;
        RECT 142.300 144.700 142.700 144.800 ;
        RECT 143.000 141.100 143.400 144.800 ;
        RECT 144.600 141.100 145.000 145.800 ;
        RECT 145.400 144.400 145.800 145.200 ;
        RECT 146.200 145.100 146.600 145.200 ;
        RECT 147.000 145.100 147.400 147.900 ;
        RECT 149.400 146.400 149.800 147.200 ;
        RECT 148.600 146.100 149.000 146.200 ;
        RECT 150.200 146.100 150.500 147.900 ;
        RECT 151.000 147.800 151.400 148.200 ;
        RECT 154.700 147.900 155.500 149.900 ;
        RECT 157.400 147.900 157.800 149.900 ;
        RECT 158.200 148.000 158.600 149.900 ;
        RECT 159.800 148.000 160.200 149.900 ;
        RECT 158.200 147.900 160.200 148.000 ;
        RECT 154.200 146.800 154.600 147.200 ;
        RECT 154.300 146.600 154.600 146.800 ;
        RECT 154.300 146.200 154.700 146.600 ;
        RECT 155.000 146.200 155.300 147.900 ;
        RECT 157.500 147.200 157.800 147.900 ;
        RECT 158.300 147.700 160.100 147.900 ;
        RECT 160.600 147.800 161.000 148.600 ;
        RECT 159.400 147.200 159.800 147.400 ;
        RECT 155.800 146.400 156.200 147.200 ;
        RECT 157.400 146.800 158.700 147.200 ;
        RECT 159.400 146.900 160.200 147.200 ;
        RECT 159.800 146.800 160.200 146.900 ;
        RECT 161.400 147.100 161.800 149.900 ;
        RECT 163.500 148.200 163.900 149.900 ;
        RECT 163.000 147.900 163.900 148.200 ;
        RECT 164.600 148.000 165.000 149.900 ;
        RECT 166.200 148.000 166.600 149.900 ;
        RECT 164.600 147.900 166.600 148.000 ;
        RECT 167.000 147.900 167.400 149.900 ;
        RECT 169.100 147.900 169.900 149.900 ;
        RECT 173.100 148.200 173.500 149.900 ;
        RECT 174.300 148.200 174.700 148.600 ;
        RECT 172.600 147.900 173.500 148.200 ;
        RECT 162.200 147.100 162.600 147.600 ;
        RECT 161.400 146.800 162.600 147.100 ;
        RECT 151.000 146.100 151.400 146.200 ;
        RECT 153.400 146.100 153.800 146.200 ;
        RECT 146.200 144.800 147.400 145.100 ;
        RECT 147.000 141.100 147.400 144.800 ;
        RECT 147.800 145.800 149.400 146.100 ;
        RECT 150.200 145.800 153.800 146.100 ;
        RECT 147.800 145.200 148.100 145.800 ;
        RECT 149.000 145.600 149.400 145.800 ;
        RECT 147.800 144.400 148.200 145.200 ;
        RECT 151.000 145.100 151.300 145.800 ;
        RECT 153.400 145.400 153.800 145.800 ;
        RECT 155.000 145.800 155.400 146.200 ;
        RECT 156.600 146.100 157.000 146.200 ;
        RECT 158.400 146.100 158.700 146.800 ;
        RECT 156.200 145.800 158.700 146.100 ;
        RECT 159.000 145.800 159.400 146.600 ;
        RECT 155.000 145.700 155.300 145.800 ;
        RECT 154.300 145.400 155.300 145.700 ;
        RECT 156.200 145.600 156.600 145.800 ;
        RECT 154.300 145.100 154.600 145.400 ;
        RECT 157.400 145.100 157.800 145.200 ;
        RECT 158.400 145.100 158.700 145.800 ;
        RECT 148.600 144.800 150.600 145.100 ;
        RECT 148.600 141.100 149.000 144.800 ;
        RECT 150.200 141.100 150.600 144.800 ;
        RECT 151.000 141.100 151.400 145.100 ;
        RECT 153.400 141.400 153.800 145.100 ;
        RECT 154.200 141.700 154.600 145.100 ;
        RECT 155.000 144.800 157.000 145.100 ;
        RECT 157.400 144.800 158.100 145.100 ;
        RECT 158.400 144.800 158.900 145.100 ;
        RECT 155.000 141.400 155.400 144.800 ;
        RECT 153.400 141.100 155.400 141.400 ;
        RECT 156.600 141.100 157.000 144.800 ;
        RECT 157.800 144.200 158.100 144.800 ;
        RECT 157.800 143.800 158.200 144.200 ;
        RECT 158.500 141.100 158.900 144.800 ;
        RECT 161.400 141.100 161.800 146.800 ;
        RECT 163.000 146.100 163.400 147.900 ;
        RECT 164.700 147.700 166.500 147.900 ;
        RECT 165.000 147.200 165.400 147.400 ;
        RECT 167.000 147.200 167.300 147.900 ;
        RECT 164.600 146.900 165.400 147.200 ;
        RECT 164.600 146.800 165.000 146.900 ;
        RECT 166.100 146.800 167.400 147.200 ;
        RECT 168.600 146.800 169.000 147.200 ;
        RECT 165.400 146.100 165.800 146.600 ;
        RECT 163.000 145.800 165.800 146.100 ;
        RECT 166.100 146.100 166.400 146.800 ;
        RECT 168.700 146.600 169.000 146.800 ;
        RECT 168.700 146.200 169.100 146.600 ;
        RECT 169.400 146.200 169.700 147.900 ;
        RECT 170.200 147.100 170.600 147.200 ;
        RECT 171.000 147.100 171.400 147.200 ;
        RECT 170.200 146.800 171.400 147.100 ;
        RECT 171.800 146.800 172.200 147.600 ;
        RECT 170.200 146.400 170.600 146.800 ;
        RECT 167.800 146.100 168.200 146.200 ;
        RECT 166.100 145.800 168.200 146.100 ;
        RECT 163.000 141.100 163.400 145.800 ;
        RECT 163.800 144.400 164.200 145.200 ;
        RECT 166.100 145.100 166.400 145.800 ;
        RECT 167.800 145.400 168.200 145.800 ;
        RECT 169.400 145.800 169.800 146.200 ;
        RECT 171.000 146.100 171.400 146.200 ;
        RECT 170.600 145.800 171.400 146.100 ;
        RECT 169.400 145.700 169.700 145.800 ;
        RECT 168.700 145.400 169.700 145.700 ;
        RECT 170.600 145.600 171.000 145.800 ;
        RECT 167.000 145.100 167.400 145.200 ;
        RECT 168.700 145.100 169.000 145.400 ;
        RECT 165.900 144.800 166.400 145.100 ;
        RECT 166.700 144.800 167.400 145.100 ;
        RECT 165.900 141.100 166.300 144.800 ;
        RECT 166.700 144.200 167.000 144.800 ;
        RECT 166.600 143.800 167.000 144.200 ;
        RECT 167.800 141.400 168.200 145.100 ;
        RECT 168.600 141.700 169.000 145.100 ;
        RECT 169.400 144.800 171.400 145.100 ;
        RECT 169.400 141.400 169.800 144.800 ;
        RECT 167.800 141.100 169.800 141.400 ;
        RECT 171.000 141.100 171.400 144.800 ;
        RECT 172.600 141.100 173.000 147.900 ;
        RECT 174.200 147.800 174.600 148.200 ;
        RECT 175.000 147.900 175.400 149.900 ;
        RECT 178.700 148.200 179.100 149.900 ;
        RECT 173.400 147.100 173.800 147.200 ;
        RECT 175.100 147.100 175.400 147.900 ;
        RECT 178.200 147.900 179.100 148.200 ;
        RECT 180.600 148.900 181.000 149.900 ;
        RECT 173.400 146.800 175.400 147.100 ;
        RECT 174.200 146.100 174.600 146.200 ;
        RECT 175.100 146.100 175.400 146.800 ;
        RECT 175.800 147.100 176.200 147.200 ;
        RECT 177.400 147.100 177.800 147.600 ;
        RECT 175.800 146.800 177.800 147.100 ;
        RECT 175.800 146.400 176.200 146.800 ;
        RECT 176.600 146.100 177.000 146.200 ;
        RECT 174.200 145.800 175.400 146.100 ;
        RECT 176.200 145.800 177.000 146.100 ;
        RECT 173.400 144.400 173.800 145.200 ;
        RECT 174.300 145.100 174.600 145.800 ;
        RECT 176.200 145.600 176.600 145.800 ;
        RECT 174.200 141.100 174.600 145.100 ;
        RECT 175.000 144.800 177.000 145.100 ;
        RECT 175.000 141.100 175.400 144.800 ;
        RECT 176.600 141.100 177.000 144.800 ;
        RECT 178.200 141.100 178.600 147.900 ;
        RECT 180.600 147.200 180.900 148.900 ;
        RECT 181.400 147.800 181.800 148.600 ;
        RECT 183.700 147.900 184.500 149.900 ;
        RECT 187.000 148.900 187.400 149.900 ;
        RECT 189.900 149.200 190.300 149.900 ;
        RECT 180.600 147.100 181.000 147.200 ;
        RECT 182.200 147.100 182.600 147.200 ;
        RECT 180.600 146.800 182.600 147.100 ;
        RECT 179.800 145.400 180.200 146.200 ;
        RECT 179.000 144.400 179.400 145.200 ;
        RECT 180.600 145.100 180.900 146.800 ;
        RECT 183.000 146.400 183.400 147.200 ;
        RECT 183.900 146.200 184.200 147.900 ;
        RECT 187.000 147.200 187.300 148.900 ;
        RECT 189.400 148.800 190.300 149.200 ;
        RECT 191.800 148.900 192.200 149.900 ;
        RECT 187.800 147.800 188.200 148.600 ;
        RECT 189.900 148.200 190.300 148.800 ;
        RECT 189.400 147.900 190.300 148.200 ;
        RECT 184.600 146.800 185.000 147.200 ;
        RECT 187.000 146.800 187.400 147.200 ;
        RECT 188.600 146.800 189.000 147.600 ;
        RECT 184.600 146.600 184.900 146.800 ;
        RECT 184.500 146.200 184.900 146.600 ;
        RECT 182.200 146.100 182.600 146.200 ;
        RECT 182.200 145.800 183.000 146.100 ;
        RECT 183.800 145.800 184.200 146.200 ;
        RECT 182.600 145.600 183.000 145.800 ;
        RECT 183.900 145.700 184.200 145.800 ;
        RECT 183.900 145.400 184.900 145.700 ;
        RECT 185.400 145.400 185.800 146.200 ;
        RECT 186.200 145.400 186.600 146.200 ;
        RECT 184.600 145.100 184.900 145.400 ;
        RECT 187.000 145.100 187.300 146.800 ;
        RECT 188.600 146.100 189.000 146.200 ;
        RECT 189.400 146.100 189.800 147.900 ;
        RECT 191.000 147.800 191.400 148.600 ;
        RECT 191.900 147.200 192.200 148.900 ;
        RECT 191.800 146.800 192.200 147.200 ;
        RECT 195.200 148.200 195.600 149.900 ;
        RECT 197.200 149.200 197.600 149.900 ;
        RECT 200.100 149.200 200.500 149.900 ;
        RECT 196.600 148.800 197.600 149.200 ;
        RECT 199.800 148.800 200.500 149.200 ;
        RECT 195.200 147.800 196.200 148.200 ;
        RECT 195.200 147.100 195.600 147.800 ;
        RECT 197.200 147.100 197.600 148.800 ;
        RECT 200.100 148.400 200.500 148.800 ;
        RECT 195.200 146.900 196.100 147.100 ;
        RECT 195.300 146.800 196.100 146.900 ;
        RECT 191.900 146.100 192.200 146.800 ;
        RECT 188.600 145.800 189.800 146.100 ;
        RECT 180.100 144.700 181.000 145.100 ;
        RECT 182.200 144.800 184.200 145.100 ;
        RECT 180.100 144.200 180.500 144.700 ;
        RECT 180.100 143.800 181.000 144.200 ;
        RECT 180.100 141.100 180.500 143.800 ;
        RECT 182.200 141.100 182.600 144.800 ;
        RECT 183.800 141.400 184.200 144.800 ;
        RECT 184.600 141.700 185.000 145.100 ;
        RECT 185.400 141.400 185.800 145.100 ;
        RECT 186.500 144.700 187.400 145.100 ;
        RECT 186.500 144.200 186.900 144.700 ;
        RECT 186.200 143.800 186.900 144.200 ;
        RECT 183.800 141.100 185.800 141.400 ;
        RECT 186.500 141.100 186.900 143.800 ;
        RECT 189.400 141.100 189.800 145.800 ;
        RECT 190.200 145.800 192.200 146.100 ;
        RECT 190.200 145.200 190.500 145.800 ;
        RECT 190.200 144.400 190.600 145.200 ;
        RECT 191.900 145.100 192.200 145.800 ;
        RECT 192.600 145.400 193.000 146.200 ;
        RECT 194.200 145.800 195.000 146.200 ;
        RECT 191.800 144.700 192.700 145.100 ;
        RECT 193.400 144.800 193.800 145.600 ;
        RECT 195.800 145.200 196.100 146.800 ;
        RECT 196.700 146.900 197.600 147.100 ;
        RECT 199.800 147.900 200.500 148.400 ;
        RECT 202.200 147.900 202.600 149.900 ;
        RECT 196.700 146.800 197.500 146.900 ;
        RECT 196.700 145.200 197.000 146.800 ;
        RECT 199.800 146.200 200.100 147.900 ;
        RECT 202.200 147.800 202.500 147.900 ;
        RECT 201.600 147.600 202.500 147.800 ;
        RECT 204.600 147.600 205.000 149.900 ;
        RECT 200.400 147.500 202.500 147.600 ;
        RECT 200.400 147.300 201.900 147.500 ;
        RECT 203.900 147.300 205.000 147.600 ;
        RECT 200.400 147.200 200.800 147.300 ;
        RECT 197.400 145.800 198.600 146.200 ;
        RECT 199.800 145.800 200.200 146.200 ;
        RECT 195.800 144.800 196.200 145.200 ;
        RECT 196.600 144.800 197.000 145.200 ;
        RECT 199.000 144.800 199.400 145.600 ;
        RECT 199.800 145.100 200.100 145.800 ;
        RECT 200.500 145.500 200.800 147.200 ;
        RECT 202.200 146.400 202.600 147.200 ;
        RECT 203.900 145.800 204.200 147.300 ;
        RECT 204.600 145.800 205.000 146.600 ;
        RECT 200.500 145.200 201.700 145.500 ;
        RECT 203.600 145.400 204.200 145.800 ;
        RECT 192.300 144.100 192.700 144.700 ;
        RECT 195.000 144.100 195.400 144.600 ;
        RECT 192.300 143.800 195.400 144.100 ;
        RECT 192.300 141.100 192.700 143.800 ;
        RECT 195.800 143.500 196.100 144.800 ;
        RECT 194.300 143.200 196.100 143.500 ;
        RECT 194.300 143.100 194.600 143.200 ;
        RECT 194.200 141.100 194.600 143.100 ;
        RECT 195.800 143.100 196.100 143.200 ;
        RECT 196.700 143.500 197.000 144.800 ;
        RECT 197.400 143.800 197.800 144.600 ;
        RECT 196.700 143.200 198.500 143.500 ;
        RECT 196.700 143.100 197.000 143.200 ;
        RECT 195.800 141.100 196.200 143.100 ;
        RECT 196.600 141.100 197.000 143.100 ;
        RECT 198.200 143.100 198.500 143.200 ;
        RECT 198.200 141.100 198.600 143.100 ;
        RECT 199.800 141.100 200.200 145.100 ;
        RECT 201.400 143.100 201.700 145.200 ;
        RECT 203.900 145.100 204.200 145.400 ;
        RECT 203.900 144.800 205.000 145.100 ;
        RECT 201.400 141.100 201.800 143.100 ;
        RECT 204.600 141.100 205.000 144.800 ;
        RECT 1.400 136.000 1.800 139.900 ;
        RECT 3.000 137.600 3.400 139.900 ;
        RECT 1.300 135.600 1.800 136.000 ;
        RECT 2.100 137.300 3.400 137.600 ;
        RECT 2.100 136.500 2.400 137.300 ;
        RECT 4.600 137.200 5.000 139.900 ;
        RECT 6.200 138.500 6.600 139.900 ;
        RECT 7.000 138.500 7.400 139.900 ;
        RECT 7.800 138.500 8.200 139.900 ;
        RECT 5.300 137.200 7.400 137.600 ;
        RECT 3.700 136.800 5.000 137.200 ;
        RECT 8.600 136.800 9.000 139.900 ;
        RECT 10.200 137.500 10.600 139.900 ;
        RECT 11.800 137.500 12.200 139.900 ;
        RECT 12.600 138.500 13.000 139.900 ;
        RECT 13.400 138.500 13.800 139.900 ;
        RECT 15.000 137.600 15.400 139.900 ;
        RECT 16.600 138.200 17.000 139.900 ;
        RECT 16.600 137.900 17.100 138.200 ;
        RECT 16.800 137.600 17.100 137.900 ;
        RECT 14.400 137.200 16.500 137.600 ;
        RECT 16.800 137.300 17.800 137.600 ;
        RECT 10.200 136.800 11.500 137.200 ;
        RECT 11.800 136.900 14.700 137.200 ;
        RECT 16.200 137.000 16.500 137.200 ;
        RECT 6.200 136.500 6.600 136.600 ;
        RECT 2.100 136.200 6.600 136.500 ;
        RECT 7.800 136.500 8.200 136.600 ;
        RECT 11.800 136.500 12.100 136.900 ;
        RECT 15.000 136.600 15.700 136.900 ;
        RECT 16.200 136.600 17.000 137.000 ;
        RECT 7.800 136.200 12.100 136.500 ;
        RECT 12.600 136.500 15.700 136.600 ;
        RECT 12.600 136.300 15.300 136.500 ;
        RECT 12.600 136.200 13.000 136.300 ;
        RECT 1.300 133.400 1.700 135.600 ;
        RECT 2.100 135.300 2.400 136.200 ;
        RECT 2.000 135.000 2.400 135.300 ;
        RECT 5.400 135.000 17.100 135.300 ;
        RECT 2.000 134.000 2.300 135.000 ;
        RECT 5.400 134.700 5.800 135.000 ;
        RECT 14.200 134.800 14.600 135.000 ;
        RECT 15.800 134.800 16.200 135.000 ;
        RECT 16.700 134.900 17.100 135.000 ;
        RECT 2.600 134.300 4.500 134.700 ;
        RECT 2.000 133.700 2.600 134.000 ;
        RECT 1.300 133.000 1.800 133.400 ;
        RECT 1.400 131.100 1.800 133.000 ;
        RECT 2.200 131.100 2.600 133.700 ;
        RECT 4.100 133.700 4.500 134.300 ;
        RECT 4.100 133.400 5.000 133.700 ;
        RECT 4.600 133.100 5.000 133.400 ;
        RECT 7.000 133.200 7.400 134.600 ;
        RECT 8.600 134.300 10.200 134.700 ;
        RECT 12.100 134.300 13.100 134.700 ;
        RECT 17.400 134.500 17.800 137.300 ;
        RECT 18.200 135.800 18.600 136.600 ;
        RECT 8.400 133.900 8.800 134.000 ;
        RECT 8.400 133.600 10.600 133.900 ;
        RECT 10.200 133.500 10.600 133.600 ;
        RECT 11.000 133.400 11.400 134.200 ;
        RECT 4.600 132.700 5.800 133.100 ;
        RECT 7.000 132.800 7.500 133.200 ;
        RECT 9.000 132.800 9.800 133.200 ;
        RECT 10.200 133.100 10.600 133.200 ;
        RECT 12.100 133.100 12.500 134.300 ;
        RECT 13.400 134.100 17.800 134.500 ;
        RECT 15.100 133.400 16.600 133.800 ;
        RECT 15.100 133.100 15.500 133.400 ;
        RECT 10.200 132.800 12.500 133.100 ;
        RECT 5.400 131.100 5.800 132.700 ;
        RECT 14.200 132.700 15.500 133.100 ;
        RECT 6.200 131.100 6.600 132.500 ;
        RECT 7.000 131.100 7.400 132.500 ;
        RECT 7.800 131.100 8.200 132.500 ;
        RECT 8.600 131.100 9.000 132.500 ;
        RECT 10.200 131.100 10.600 132.500 ;
        RECT 11.800 131.100 12.200 132.500 ;
        RECT 12.600 131.100 13.000 132.500 ;
        RECT 13.400 131.100 13.800 132.500 ;
        RECT 14.200 131.100 14.600 132.700 ;
        RECT 17.400 131.100 17.800 134.100 ;
        RECT 19.000 133.100 19.400 139.900 ;
        RECT 21.400 136.000 21.800 139.900 ;
        RECT 23.000 137.600 23.400 139.900 ;
        RECT 21.300 135.600 21.800 136.000 ;
        RECT 22.100 137.300 23.400 137.600 ;
        RECT 22.100 136.500 22.400 137.300 ;
        RECT 24.600 137.200 25.000 139.900 ;
        RECT 26.200 138.500 26.600 139.900 ;
        RECT 27.000 138.500 27.400 139.900 ;
        RECT 27.800 138.500 28.200 139.900 ;
        RECT 25.300 137.200 27.400 137.600 ;
        RECT 23.700 136.800 25.000 137.200 ;
        RECT 28.600 136.800 29.000 139.900 ;
        RECT 30.200 137.500 30.600 139.900 ;
        RECT 31.800 137.500 32.200 139.900 ;
        RECT 32.600 138.500 33.000 139.900 ;
        RECT 33.400 138.500 33.800 139.900 ;
        RECT 35.000 137.600 35.400 139.900 ;
        RECT 36.600 138.200 37.000 139.900 ;
        RECT 36.600 137.900 37.100 138.200 ;
        RECT 36.800 137.600 37.100 137.900 ;
        RECT 34.400 137.200 36.500 137.600 ;
        RECT 36.800 137.300 37.800 137.600 ;
        RECT 30.200 136.800 31.500 137.200 ;
        RECT 31.800 136.900 34.700 137.200 ;
        RECT 36.200 137.000 36.500 137.200 ;
        RECT 26.200 136.500 26.600 136.600 ;
        RECT 22.100 136.200 26.600 136.500 ;
        RECT 27.800 136.500 28.200 136.600 ;
        RECT 31.800 136.500 32.100 136.900 ;
        RECT 35.000 136.600 35.700 136.900 ;
        RECT 36.200 136.600 37.000 137.000 ;
        RECT 27.800 136.200 32.100 136.500 ;
        RECT 32.600 136.500 35.700 136.600 ;
        RECT 32.600 136.300 35.300 136.500 ;
        RECT 32.600 136.200 33.000 136.300 ;
        RECT 19.800 133.400 20.200 134.200 ;
        RECT 21.300 133.400 21.700 135.600 ;
        RECT 22.100 135.300 22.400 136.200 ;
        RECT 22.000 135.000 22.400 135.300 ;
        RECT 25.400 135.000 37.100 135.300 ;
        RECT 22.000 134.000 22.300 135.000 ;
        RECT 25.400 134.700 25.800 135.000 ;
        RECT 34.200 134.800 34.600 135.000 ;
        RECT 36.700 134.900 37.100 135.000 ;
        RECT 22.600 134.300 24.500 134.700 ;
        RECT 22.000 133.700 22.600 134.000 ;
        RECT 18.500 132.800 19.400 133.100 ;
        RECT 21.300 133.000 21.800 133.400 ;
        RECT 18.500 131.100 18.900 132.800 ;
        RECT 21.400 131.100 21.800 133.000 ;
        RECT 22.200 131.100 22.600 133.700 ;
        RECT 24.100 133.700 24.500 134.300 ;
        RECT 24.100 133.400 25.000 133.700 ;
        RECT 24.600 133.100 25.000 133.400 ;
        RECT 27.000 133.200 27.400 134.600 ;
        RECT 28.600 134.300 30.200 134.700 ;
        RECT 32.100 134.300 33.100 134.700 ;
        RECT 37.400 134.500 37.800 137.300 ;
        RECT 39.500 136.200 39.900 139.900 ;
        RECT 40.200 136.800 40.600 137.200 ;
        RECT 40.300 136.200 40.600 136.800 ;
        RECT 41.400 136.200 41.800 139.900 ;
        RECT 43.000 136.200 43.400 139.900 ;
        RECT 39.500 135.900 40.000 136.200 ;
        RECT 40.300 135.900 41.000 136.200 ;
        RECT 41.400 135.900 43.400 136.200 ;
        RECT 43.800 135.900 44.200 139.900 ;
        RECT 45.000 136.800 45.400 137.200 ;
        RECT 45.000 136.200 45.300 136.800 ;
        RECT 45.700 136.200 46.100 139.900 ;
        RECT 44.600 135.900 45.300 136.200 ;
        RECT 45.600 135.900 46.100 136.200 ;
        RECT 47.800 135.900 48.200 139.900 ;
        RECT 48.600 136.200 49.000 139.900 ;
        RECT 50.200 136.200 50.600 139.900 ;
        RECT 48.600 135.900 50.600 136.200 ;
        RECT 28.400 133.900 28.800 134.000 ;
        RECT 28.400 133.600 30.600 133.900 ;
        RECT 30.200 133.500 30.600 133.600 ;
        RECT 31.000 133.400 31.400 134.200 ;
        RECT 24.600 132.700 25.800 133.100 ;
        RECT 27.000 132.800 27.500 133.200 ;
        RECT 29.000 132.800 29.800 133.200 ;
        RECT 30.200 133.100 30.600 133.200 ;
        RECT 32.100 133.100 32.500 134.300 ;
        RECT 33.400 134.100 37.800 134.500 ;
        RECT 39.000 134.400 39.400 135.200 ;
        RECT 39.700 134.200 40.000 135.900 ;
        RECT 40.600 135.800 41.000 135.900 ;
        RECT 41.800 135.200 42.200 135.400 ;
        RECT 43.800 135.200 44.100 135.900 ;
        RECT 44.600 135.800 45.000 135.900 ;
        RECT 41.400 134.900 42.200 135.200 ;
        RECT 43.000 134.900 44.200 135.200 ;
        RECT 41.400 134.800 41.800 134.900 ;
        RECT 35.100 133.400 36.600 133.800 ;
        RECT 35.100 133.100 35.500 133.400 ;
        RECT 30.200 132.800 32.500 133.100 ;
        RECT 25.400 131.100 25.800 132.700 ;
        RECT 34.200 132.700 35.500 133.100 ;
        RECT 26.200 131.100 26.600 132.500 ;
        RECT 27.000 131.100 27.400 132.500 ;
        RECT 27.800 131.100 28.200 132.500 ;
        RECT 28.600 131.100 29.000 132.500 ;
        RECT 30.200 131.100 30.600 132.500 ;
        RECT 31.800 131.100 32.200 132.500 ;
        RECT 32.600 131.100 33.000 132.500 ;
        RECT 33.400 131.100 33.800 132.500 ;
        RECT 34.200 131.100 34.600 132.700 ;
        RECT 37.400 131.100 37.800 134.100 ;
        RECT 38.200 134.100 38.600 134.200 ;
        RECT 38.200 133.800 39.000 134.100 ;
        RECT 39.700 133.800 41.000 134.200 ;
        RECT 42.200 133.800 42.600 134.600 ;
        RECT 38.600 133.600 39.000 133.800 ;
        RECT 38.300 133.100 40.100 133.300 ;
        RECT 40.600 133.100 40.900 133.800 ;
        RECT 43.000 133.100 43.300 134.900 ;
        RECT 43.800 134.800 44.200 134.900 ;
        RECT 45.600 134.200 45.900 135.900 ;
        RECT 47.900 135.200 48.200 135.900 ;
        RECT 52.600 135.700 53.000 139.900 ;
        RECT 54.800 138.200 55.200 139.900 ;
        RECT 54.200 137.900 55.200 138.200 ;
        RECT 57.000 137.900 57.400 139.900 ;
        RECT 59.100 137.900 59.700 139.900 ;
        RECT 54.200 137.500 54.600 137.900 ;
        RECT 57.000 137.600 57.300 137.900 ;
        RECT 55.900 137.300 57.700 137.600 ;
        RECT 59.000 137.500 59.400 137.900 ;
        RECT 55.900 137.200 56.300 137.300 ;
        RECT 57.300 137.200 57.700 137.300 ;
        RECT 61.400 137.100 61.800 139.900 ;
        RECT 62.200 137.100 62.600 137.200 ;
        RECT 54.200 136.500 54.600 136.600 ;
        RECT 56.500 136.500 56.900 136.600 ;
        RECT 54.200 136.200 56.900 136.500 ;
        RECT 57.200 136.500 58.300 136.800 ;
        RECT 57.200 135.900 57.500 136.500 ;
        RECT 57.900 136.400 58.300 136.500 ;
        RECT 59.100 136.600 59.800 137.000 ;
        RECT 61.400 136.800 62.600 137.100 ;
        RECT 59.100 136.100 59.400 136.600 ;
        RECT 55.100 135.700 57.500 135.900 ;
        RECT 52.600 135.600 57.500 135.700 ;
        RECT 58.200 135.800 59.400 136.100 ;
        RECT 52.600 135.500 55.500 135.600 ;
        RECT 52.600 135.400 55.400 135.500 ;
        RECT 49.800 135.200 50.200 135.400 ;
        RECT 46.200 134.400 46.600 135.200 ;
        RECT 47.800 134.900 49.000 135.200 ;
        RECT 49.800 134.900 50.600 135.200 ;
        RECT 55.800 135.100 56.200 135.200 ;
        RECT 47.800 134.800 48.200 134.900 ;
        RECT 44.600 133.800 45.900 134.200 ;
        RECT 47.000 134.100 47.400 134.200 ;
        RECT 46.600 133.800 47.400 134.100 ;
        RECT 38.200 133.000 40.200 133.100 ;
        RECT 38.200 131.100 38.600 133.000 ;
        RECT 39.800 131.100 40.200 133.000 ;
        RECT 40.600 131.100 41.000 133.100 ;
        RECT 43.000 131.100 43.400 133.100 ;
        RECT 43.800 132.800 44.200 133.200 ;
        RECT 44.700 133.100 45.000 133.800 ;
        RECT 46.600 133.600 47.000 133.800 ;
        RECT 45.500 133.100 47.300 133.300 ;
        RECT 43.700 132.400 44.100 132.800 ;
        RECT 44.600 131.100 45.000 133.100 ;
        RECT 45.400 133.000 47.400 133.100 ;
        RECT 45.400 131.100 45.800 133.000 ;
        RECT 47.000 131.100 47.400 133.000 ;
        RECT 47.800 132.800 48.200 133.200 ;
        RECT 48.700 133.100 49.000 134.900 ;
        RECT 50.200 134.800 50.600 134.900 ;
        RECT 53.700 134.800 56.200 135.100 ;
        RECT 53.700 134.700 54.100 134.800 ;
        RECT 49.400 134.100 49.800 134.600 ;
        RECT 54.500 134.200 54.900 134.300 ;
        RECT 58.200 134.200 58.500 135.800 ;
        RECT 61.400 135.600 61.800 136.800 ;
        RECT 59.700 135.300 61.800 135.600 ;
        RECT 59.700 135.200 60.100 135.300 ;
        RECT 60.500 134.900 60.900 135.000 ;
        RECT 59.000 134.600 60.900 134.900 ;
        RECT 59.000 134.500 59.400 134.600 ;
        RECT 51.800 134.100 52.200 134.200 ;
        RECT 49.400 133.800 52.200 134.100 ;
        RECT 53.000 133.900 58.500 134.200 ;
        RECT 53.000 133.800 53.800 133.900 ;
        RECT 47.900 132.400 48.300 132.800 ;
        RECT 48.600 131.100 49.000 133.100 ;
        RECT 52.600 131.100 53.000 133.500 ;
        RECT 55.100 133.200 55.400 133.900 ;
        RECT 57.900 133.800 58.300 133.900 ;
        RECT 61.400 133.600 61.800 135.300 ;
        RECT 63.000 135.100 63.400 139.900 ;
        RECT 65.000 136.800 65.400 137.200 ;
        RECT 63.800 135.800 64.200 136.600 ;
        RECT 65.000 136.200 65.300 136.800 ;
        RECT 65.700 136.200 66.100 139.900 ;
        RECT 64.600 135.900 65.300 136.200 ;
        RECT 65.600 135.900 66.100 136.200 ;
        RECT 69.100 136.200 69.500 139.900 ;
        RECT 69.800 136.800 70.200 137.200 ;
        RECT 69.900 136.200 70.200 136.800 ;
        RECT 69.100 135.900 69.600 136.200 ;
        RECT 69.900 135.900 70.600 136.200 ;
        RECT 64.600 135.800 65.000 135.900 ;
        RECT 64.600 135.100 64.900 135.800 ;
        RECT 65.600 135.200 65.900 135.900 ;
        RECT 63.000 134.800 64.900 135.100 ;
        RECT 65.400 134.800 65.900 135.200 ;
        RECT 59.900 133.300 61.800 133.600 ;
        RECT 62.200 133.400 62.600 134.200 ;
        RECT 59.900 133.200 60.300 133.300 ;
        RECT 54.200 132.100 54.600 132.500 ;
        RECT 55.000 132.400 55.400 133.200 ;
        RECT 55.900 132.700 56.300 132.800 ;
        RECT 55.900 132.400 57.300 132.700 ;
        RECT 57.000 132.100 57.300 132.400 ;
        RECT 59.000 132.100 59.400 132.500 ;
        RECT 54.200 131.800 55.200 132.100 ;
        RECT 54.800 131.100 55.200 131.800 ;
        RECT 57.000 131.100 57.400 132.100 ;
        RECT 59.000 131.800 59.700 132.100 ;
        RECT 59.100 131.100 59.700 131.800 ;
        RECT 61.400 131.100 61.800 133.300 ;
        RECT 63.000 133.100 63.400 134.800 ;
        RECT 65.600 134.200 65.900 134.800 ;
        RECT 66.200 134.400 66.600 135.200 ;
        RECT 67.000 135.100 67.400 135.200 ;
        RECT 68.600 135.100 69.000 135.200 ;
        RECT 67.000 134.800 69.000 135.100 ;
        RECT 68.600 134.400 69.000 134.800 ;
        RECT 69.300 134.200 69.600 135.900 ;
        RECT 70.200 135.800 70.600 135.900 ;
        RECT 71.000 135.800 71.400 136.600 ;
        RECT 64.600 133.800 65.900 134.200 ;
        RECT 67.000 134.100 67.400 134.200 ;
        RECT 66.600 133.800 67.400 134.100 ;
        RECT 67.800 134.100 68.200 134.200 ;
        RECT 67.800 133.800 68.600 134.100 ;
        RECT 69.300 133.800 70.600 134.200 ;
        RECT 64.700 133.100 65.000 133.800 ;
        RECT 66.600 133.600 67.000 133.800 ;
        RECT 68.200 133.600 68.600 133.800 ;
        RECT 65.500 133.100 67.300 133.300 ;
        RECT 67.900 133.100 69.700 133.300 ;
        RECT 70.200 133.100 70.500 133.800 ;
        RECT 71.800 133.100 72.200 139.900 ;
        RECT 73.400 136.200 73.800 139.900 ;
        RECT 75.000 136.200 75.400 139.900 ;
        RECT 73.400 135.900 75.400 136.200 ;
        RECT 75.800 135.900 76.200 139.900 ;
        RECT 73.800 135.200 74.200 135.400 ;
        RECT 75.800 135.200 76.100 135.900 ;
        RECT 73.400 134.900 74.200 135.200 ;
        RECT 75.000 134.900 76.200 135.200 ;
        RECT 73.400 134.800 73.800 134.900 ;
        RECT 72.600 133.400 73.000 134.200 ;
        RECT 74.200 133.800 74.600 134.600 ;
        RECT 63.000 132.800 63.900 133.100 ;
        RECT 63.500 131.100 63.900 132.800 ;
        RECT 64.600 131.100 65.000 133.100 ;
        RECT 65.400 133.000 67.400 133.100 ;
        RECT 65.400 131.100 65.800 133.000 ;
        RECT 67.000 131.100 67.400 133.000 ;
        RECT 67.800 133.000 69.800 133.100 ;
        RECT 67.800 131.100 68.200 133.000 ;
        RECT 69.400 131.100 69.800 133.000 ;
        RECT 70.200 131.100 70.600 133.100 ;
        RECT 71.300 132.800 72.200 133.100 ;
        RECT 75.000 133.100 75.300 134.900 ;
        RECT 75.800 134.800 76.200 134.900 ;
        RECT 77.400 135.100 77.800 139.900 ;
        RECT 79.400 136.800 79.800 137.200 ;
        RECT 78.200 135.800 78.600 136.600 ;
        RECT 79.400 136.200 79.700 136.800 ;
        RECT 80.100 136.200 80.500 139.900 ;
        RECT 79.000 135.900 79.700 136.200 ;
        RECT 80.000 135.900 80.500 136.200 ;
        RECT 79.000 135.800 79.400 135.900 ;
        RECT 79.000 135.100 79.300 135.800 ;
        RECT 80.000 135.200 80.300 135.900 ;
        RECT 82.200 135.600 82.600 139.900 ;
        RECT 84.300 137.900 84.900 139.900 ;
        RECT 86.600 137.900 87.000 139.900 ;
        RECT 88.800 138.200 89.200 139.900 ;
        RECT 88.800 137.900 89.800 138.200 ;
        RECT 84.600 137.500 85.000 137.900 ;
        RECT 86.700 137.600 87.000 137.900 ;
        RECT 86.300 137.300 88.100 137.600 ;
        RECT 89.400 137.500 89.800 137.900 ;
        RECT 86.300 137.200 86.700 137.300 ;
        RECT 87.700 137.200 88.100 137.300 ;
        RECT 84.200 136.600 84.900 137.000 ;
        RECT 84.600 136.100 84.900 136.600 ;
        RECT 85.700 136.500 86.800 136.800 ;
        RECT 85.700 136.400 86.100 136.500 ;
        RECT 84.600 135.800 85.800 136.100 ;
        RECT 82.200 135.300 84.300 135.600 ;
        RECT 77.400 134.800 79.300 135.100 ;
        RECT 79.800 134.800 80.300 135.200 ;
        RECT 76.600 133.400 77.000 134.200 ;
        RECT 71.300 132.200 71.700 132.800 ;
        RECT 71.300 131.800 72.200 132.200 ;
        RECT 71.300 131.100 71.700 131.800 ;
        RECT 75.000 131.100 75.400 133.100 ;
        RECT 75.800 132.800 76.200 133.200 ;
        RECT 77.400 133.100 77.800 134.800 ;
        RECT 80.000 134.200 80.300 134.800 ;
        RECT 80.600 134.400 81.000 135.200 ;
        RECT 79.000 133.800 80.300 134.200 ;
        RECT 81.400 134.100 81.800 134.200 ;
        RECT 81.000 133.800 81.800 134.100 ;
        RECT 79.100 133.100 79.400 133.800 ;
        RECT 81.000 133.600 81.400 133.800 ;
        RECT 82.200 133.600 82.600 135.300 ;
        RECT 83.900 135.200 84.300 135.300 ;
        RECT 83.100 134.900 83.500 135.000 ;
        RECT 83.100 134.600 85.000 134.900 ;
        RECT 84.600 134.500 85.000 134.600 ;
        RECT 85.500 134.200 85.800 135.800 ;
        RECT 86.500 135.900 86.800 136.500 ;
        RECT 87.100 136.500 87.500 136.600 ;
        RECT 89.400 136.500 89.800 136.600 ;
        RECT 87.100 136.200 89.800 136.500 ;
        RECT 86.500 135.700 88.900 135.900 ;
        RECT 91.000 135.700 91.400 139.900 ;
        RECT 86.500 135.600 91.400 135.700 ;
        RECT 88.500 135.500 91.400 135.600 ;
        RECT 88.600 135.400 91.400 135.500 ;
        RECT 87.800 135.100 88.200 135.200 ;
        RECT 92.600 135.100 93.000 139.900 ;
        RECT 94.600 136.800 95.000 137.200 ;
        RECT 93.400 135.800 93.800 136.600 ;
        RECT 94.600 136.200 94.900 136.800 ;
        RECT 95.300 136.200 95.700 139.900 ;
        RECT 98.200 136.400 98.600 139.900 ;
        RECT 94.200 135.900 94.900 136.200 ;
        RECT 95.200 135.900 95.700 136.200 ;
        RECT 98.100 135.900 98.600 136.400 ;
        RECT 99.800 136.200 100.200 139.900 ;
        RECT 98.900 135.900 100.200 136.200 ;
        RECT 102.200 136.200 102.600 139.900 ;
        RECT 103.800 136.400 104.200 139.900 ;
        RECT 105.400 137.500 105.800 139.500 ;
        RECT 102.200 135.900 103.500 136.200 ;
        RECT 103.800 135.900 104.300 136.400 ;
        RECT 94.200 135.800 94.600 135.900 ;
        RECT 94.200 135.100 94.500 135.800 ;
        RECT 87.800 134.800 90.300 135.100 ;
        RECT 88.600 134.700 89.000 134.800 ;
        RECT 89.900 134.700 90.300 134.800 ;
        RECT 92.600 134.800 94.500 135.100 ;
        RECT 89.100 134.200 89.500 134.300 ;
        RECT 85.500 133.900 91.000 134.200 ;
        RECT 85.700 133.800 86.100 133.900 ;
        RECT 87.000 133.800 87.400 133.900 ;
        RECT 82.200 133.300 84.100 133.600 ;
        RECT 79.900 133.100 81.700 133.300 ;
        RECT 77.400 132.800 78.300 133.100 ;
        RECT 75.700 132.400 76.100 132.800 ;
        RECT 77.900 131.100 78.300 132.800 ;
        RECT 79.000 131.100 79.400 133.100 ;
        RECT 79.800 133.000 81.800 133.100 ;
        RECT 79.800 131.100 80.200 133.000 ;
        RECT 81.400 131.100 81.800 133.000 ;
        RECT 82.200 131.100 82.600 133.300 ;
        RECT 83.700 133.200 84.100 133.300 ;
        RECT 88.600 132.800 88.900 133.900 ;
        RECT 90.200 133.800 91.000 133.900 ;
        RECT 87.700 132.700 88.100 132.800 ;
        RECT 84.600 132.100 85.000 132.500 ;
        RECT 86.700 132.400 88.100 132.700 ;
        RECT 88.600 132.400 89.000 132.800 ;
        RECT 86.700 132.100 87.000 132.400 ;
        RECT 89.400 132.100 89.800 132.500 ;
        RECT 84.300 131.800 85.000 132.100 ;
        RECT 84.300 131.100 84.900 131.800 ;
        RECT 86.600 131.100 87.000 132.100 ;
        RECT 88.800 131.800 89.800 132.100 ;
        RECT 88.800 131.100 89.200 131.800 ;
        RECT 91.000 131.100 91.400 133.500 ;
        RECT 91.800 133.400 92.200 134.200 ;
        RECT 92.600 133.100 93.000 134.800 ;
        RECT 95.200 134.200 95.500 135.900 ;
        RECT 95.800 134.400 96.200 135.200 ;
        RECT 98.100 134.200 98.400 135.900 ;
        RECT 98.900 134.900 99.200 135.900 ;
        RECT 98.700 134.500 99.200 134.900 ;
        RECT 94.200 133.800 95.500 134.200 ;
        RECT 96.600 134.100 97.000 134.200 ;
        RECT 96.200 133.800 97.000 134.100 ;
        RECT 98.100 133.800 98.600 134.200 ;
        RECT 94.300 133.100 94.600 133.800 ;
        RECT 96.200 133.600 96.600 133.800 ;
        RECT 95.100 133.100 96.900 133.300 ;
        RECT 98.100 133.200 98.400 133.800 ;
        RECT 98.900 133.700 99.200 134.500 ;
        RECT 99.700 135.100 100.200 135.200 ;
        RECT 102.200 135.100 102.700 135.200 ;
        RECT 99.700 134.800 102.700 135.100 ;
        RECT 99.700 134.400 100.100 134.800 ;
        RECT 102.300 134.400 102.700 134.800 ;
        RECT 103.200 134.900 103.500 135.900 ;
        RECT 103.200 134.500 103.700 134.900 ;
        RECT 103.200 133.700 103.500 134.500 ;
        RECT 104.000 134.200 104.300 135.900 ;
        RECT 105.400 135.800 105.700 137.500 ;
        RECT 107.500 136.400 107.900 139.900 ;
        RECT 107.500 136.100 108.300 136.400 ;
        RECT 105.400 135.500 107.300 135.800 ;
        RECT 105.400 134.400 105.800 135.200 ;
        RECT 106.200 134.400 106.600 135.200 ;
        RECT 107.000 134.500 107.300 135.500 ;
        RECT 103.800 134.100 104.300 134.200 ;
        RECT 104.600 134.100 105.000 134.200 ;
        RECT 103.800 133.800 105.000 134.100 ;
        RECT 107.000 134.100 107.700 134.500 ;
        RECT 108.000 134.200 108.300 136.100 ;
        RECT 111.500 136.200 111.900 139.900 ;
        RECT 112.200 136.800 112.600 137.200 ;
        RECT 112.300 136.200 112.600 136.800 ;
        RECT 111.500 135.900 112.000 136.200 ;
        RECT 112.300 135.900 113.000 136.200 ;
        RECT 108.600 134.800 109.000 135.600 ;
        RECT 111.000 134.400 111.400 135.200 ;
        RECT 111.700 134.200 112.000 135.900 ;
        RECT 112.600 135.800 113.000 135.900 ;
        RECT 113.400 135.800 113.800 136.600 ;
        RECT 112.600 135.100 112.900 135.800 ;
        RECT 114.200 135.100 114.600 139.900 ;
        RECT 112.600 134.800 114.600 135.100 ;
        RECT 107.000 133.900 107.500 134.100 ;
        RECT 98.900 133.400 100.200 133.700 ;
        RECT 92.600 132.800 93.500 133.100 ;
        RECT 93.100 131.100 93.500 132.800 ;
        RECT 94.200 131.100 94.600 133.100 ;
        RECT 95.000 133.000 97.000 133.100 ;
        RECT 95.000 131.100 95.400 133.000 ;
        RECT 96.600 131.100 97.000 133.000 ;
        RECT 98.100 132.800 98.600 133.200 ;
        RECT 98.200 131.100 98.600 132.800 ;
        RECT 99.800 131.100 100.200 133.400 ;
        RECT 102.200 133.400 103.500 133.700 ;
        RECT 102.200 131.100 102.600 133.400 ;
        RECT 104.000 133.100 104.300 133.800 ;
        RECT 103.800 132.800 104.300 133.100 ;
        RECT 105.400 133.600 107.500 133.900 ;
        RECT 108.000 133.800 109.000 134.200 ;
        RECT 110.200 134.100 110.600 134.200 ;
        RECT 110.200 133.800 111.000 134.100 ;
        RECT 111.700 133.800 113.000 134.200 ;
        RECT 103.800 131.100 104.200 132.800 ;
        RECT 105.400 132.500 105.700 133.600 ;
        RECT 108.000 133.500 108.300 133.800 ;
        RECT 110.600 133.600 111.000 133.800 ;
        RECT 107.900 133.300 108.300 133.500 ;
        RECT 107.500 133.000 108.300 133.300 ;
        RECT 110.300 133.100 112.100 133.300 ;
        RECT 112.600 133.100 112.900 133.800 ;
        RECT 114.200 133.100 114.600 134.800 ;
        RECT 115.800 135.600 116.200 139.900 ;
        RECT 117.900 137.900 118.500 139.900 ;
        RECT 120.200 137.900 120.600 139.900 ;
        RECT 122.400 138.200 122.800 139.900 ;
        RECT 122.400 137.900 123.400 138.200 ;
        RECT 118.200 137.500 118.600 137.900 ;
        RECT 120.300 137.600 120.600 137.900 ;
        RECT 119.900 137.300 121.700 137.600 ;
        RECT 123.000 137.500 123.400 137.900 ;
        RECT 119.900 137.200 120.300 137.300 ;
        RECT 121.300 137.200 121.700 137.300 ;
        RECT 117.800 136.600 118.500 137.000 ;
        RECT 118.200 136.100 118.500 136.600 ;
        RECT 119.300 136.500 120.400 136.800 ;
        RECT 119.300 136.400 119.700 136.500 ;
        RECT 118.200 135.800 119.400 136.100 ;
        RECT 115.800 135.300 117.900 135.600 ;
        RECT 115.000 133.400 115.400 134.200 ;
        RECT 115.800 133.600 116.200 135.300 ;
        RECT 117.500 135.200 117.900 135.300 ;
        RECT 119.100 135.200 119.400 135.800 ;
        RECT 120.100 135.900 120.400 136.500 ;
        RECT 120.700 136.500 121.100 136.600 ;
        RECT 123.000 136.500 123.400 136.600 ;
        RECT 120.700 136.200 123.400 136.500 ;
        RECT 120.100 135.700 122.500 135.900 ;
        RECT 124.600 135.700 125.000 139.900 ;
        RECT 125.400 135.800 125.800 136.600 ;
        RECT 120.100 135.600 125.000 135.700 ;
        RECT 122.100 135.500 125.000 135.600 ;
        RECT 122.200 135.400 125.000 135.500 ;
        RECT 116.700 134.900 117.100 135.000 ;
        RECT 116.700 134.600 118.600 134.900 ;
        RECT 119.000 134.800 119.400 135.200 ;
        RECT 121.400 135.100 121.800 135.200 ;
        RECT 121.400 134.800 123.900 135.100 ;
        RECT 118.200 134.500 118.600 134.600 ;
        RECT 119.100 134.200 119.400 134.800 ;
        RECT 122.200 134.700 122.600 134.800 ;
        RECT 123.500 134.700 123.900 134.800 ;
        RECT 122.700 134.200 123.100 134.300 ;
        RECT 119.100 133.900 124.600 134.200 ;
        RECT 119.300 133.800 119.700 133.900 ;
        RECT 110.200 133.000 112.200 133.100 ;
        RECT 105.400 131.500 105.800 132.500 ;
        RECT 107.500 132.200 107.900 133.000 ;
        RECT 107.000 131.800 107.900 132.200 ;
        RECT 107.500 131.500 107.900 131.800 ;
        RECT 110.200 131.100 110.600 133.000 ;
        RECT 111.800 131.100 112.200 133.000 ;
        RECT 112.600 131.100 113.000 133.100 ;
        RECT 113.700 132.800 114.600 133.100 ;
        RECT 115.800 133.300 117.700 133.600 ;
        RECT 113.700 131.100 114.100 132.800 ;
        RECT 115.800 131.100 116.200 133.300 ;
        RECT 117.300 133.200 117.700 133.300 ;
        RECT 122.200 132.800 122.500 133.900 ;
        RECT 123.800 133.800 124.600 133.900 ;
        RECT 121.300 132.700 121.700 132.800 ;
        RECT 118.200 132.100 118.600 132.500 ;
        RECT 120.300 132.400 121.700 132.700 ;
        RECT 122.200 132.400 122.600 132.800 ;
        RECT 120.300 132.100 120.600 132.400 ;
        RECT 123.000 132.100 123.400 132.500 ;
        RECT 117.900 131.800 118.600 132.100 ;
        RECT 117.900 131.100 118.500 131.800 ;
        RECT 120.200 131.100 120.600 132.100 ;
        RECT 122.400 131.800 123.400 132.100 ;
        RECT 122.400 131.100 122.800 131.800 ;
        RECT 124.600 131.100 125.000 133.500 ;
        RECT 126.200 133.100 126.600 139.900 ;
        RECT 127.000 134.100 127.400 134.200 ;
        RECT 127.800 134.100 128.200 134.200 ;
        RECT 127.000 133.800 128.200 134.100 ;
        RECT 127.000 133.400 127.400 133.800 ;
        RECT 127.800 133.400 128.200 133.800 ;
        RECT 125.700 132.800 126.600 133.100 ;
        RECT 128.600 133.100 129.000 139.900 ;
        RECT 129.400 135.800 129.800 136.600 ;
        RECT 131.500 136.300 131.900 139.900 ;
        RECT 133.900 136.300 134.300 139.900 ;
        RECT 136.300 136.300 136.700 139.900 ;
        RECT 131.000 135.900 131.900 136.300 ;
        RECT 133.400 135.900 134.300 136.300 ;
        RECT 135.800 135.900 136.700 136.300 ;
        RECT 137.400 135.900 137.800 139.900 ;
        RECT 138.200 136.200 138.600 139.900 ;
        RECT 139.800 136.200 140.200 139.900 ;
        RECT 141.400 136.400 141.800 139.900 ;
        RECT 138.200 135.900 140.200 136.200 ;
        RECT 141.300 135.900 141.800 136.400 ;
        RECT 143.000 136.200 143.400 139.900 ;
        RECT 142.100 135.900 143.400 136.200 ;
        RECT 143.800 136.200 144.200 139.900 ;
        RECT 145.400 136.400 145.800 139.900 ;
        RECT 143.800 135.900 145.100 136.200 ;
        RECT 145.400 135.900 145.900 136.400 ;
        RECT 147.000 136.200 147.400 139.900 ;
        RECT 148.600 136.400 149.000 139.900 ;
        RECT 147.000 135.900 148.300 136.200 ;
        RECT 130.200 135.100 130.600 135.200 ;
        RECT 131.100 135.100 131.400 135.900 ;
        RECT 130.200 134.800 131.400 135.100 ;
        RECT 131.800 134.800 132.200 135.600 ;
        RECT 131.100 134.200 131.400 134.800 ;
        RECT 133.500 134.200 133.800 135.900 ;
        RECT 134.200 134.800 134.600 135.600 ;
        RECT 135.900 134.200 136.200 135.900 ;
        RECT 136.600 134.800 137.000 135.600 ;
        RECT 137.500 135.200 137.800 135.900 ;
        RECT 139.400 135.200 139.800 135.400 ;
        RECT 137.400 134.900 138.600 135.200 ;
        RECT 139.400 134.900 140.200 135.200 ;
        RECT 137.400 134.800 137.800 134.900 ;
        RECT 131.000 133.800 131.400 134.200 ;
        RECT 133.400 133.800 133.800 134.200 ;
        RECT 130.200 133.100 130.600 133.200 ;
        RECT 128.600 132.800 130.600 133.100 ;
        RECT 125.700 131.100 126.100 132.800 ;
        RECT 129.100 131.100 129.500 132.800 ;
        RECT 130.200 132.400 130.600 132.800 ;
        RECT 131.100 132.100 131.400 133.800 ;
        RECT 132.600 132.400 133.000 133.200 ;
        RECT 133.500 133.100 133.800 133.800 ;
        RECT 134.200 133.800 134.600 134.200 ;
        RECT 135.800 133.800 136.200 134.200 ;
        RECT 134.200 133.100 134.500 133.800 ;
        RECT 133.400 132.800 134.500 133.100 ;
        RECT 133.500 132.100 133.800 132.800 ;
        RECT 135.000 132.400 135.400 133.200 ;
        RECT 135.900 133.100 136.200 133.800 ;
        RECT 137.400 133.100 137.800 133.200 ;
        RECT 138.300 133.100 138.600 134.900 ;
        RECT 139.800 134.800 140.200 134.900 ;
        RECT 139.000 133.800 139.400 134.600 ;
        RECT 141.300 134.200 141.600 135.900 ;
        RECT 142.100 134.900 142.400 135.900 ;
        RECT 141.900 134.500 142.400 134.900 ;
        RECT 141.300 133.800 141.800 134.200 ;
        RECT 135.800 132.800 137.800 133.100 ;
        RECT 135.900 132.100 136.200 132.800 ;
        RECT 137.500 132.400 137.900 132.800 ;
        RECT 131.000 131.100 131.400 132.100 ;
        RECT 133.400 131.100 133.800 132.100 ;
        RECT 135.800 131.100 136.200 132.100 ;
        RECT 138.200 131.100 138.600 133.100 ;
        RECT 141.300 133.100 141.600 133.800 ;
        RECT 142.100 133.700 142.400 134.500 ;
        RECT 142.900 134.800 143.400 135.200 ;
        RECT 143.800 134.800 144.300 135.200 ;
        RECT 142.900 134.400 143.300 134.800 ;
        RECT 143.900 134.400 144.300 134.800 ;
        RECT 144.800 134.900 145.100 135.900 ;
        RECT 144.800 134.500 145.300 134.900 ;
        RECT 144.800 133.700 145.100 134.500 ;
        RECT 145.600 134.200 145.900 135.900 ;
        RECT 147.000 135.100 147.500 135.200 ;
        RECT 145.400 133.800 145.900 134.200 ;
        RECT 146.200 134.800 147.500 135.100 ;
        RECT 146.200 134.200 146.500 134.800 ;
        RECT 147.100 134.400 147.500 134.800 ;
        RECT 148.000 134.900 148.300 135.900 ;
        RECT 148.600 135.800 149.100 136.400 ;
        RECT 148.000 134.500 148.500 134.900 ;
        RECT 146.200 133.800 146.600 134.200 ;
        RECT 142.100 133.400 143.400 133.700 ;
        RECT 141.300 132.800 141.800 133.100 ;
        RECT 141.400 131.100 141.800 132.800 ;
        RECT 143.000 131.100 143.400 133.400 ;
        RECT 143.800 133.400 145.100 133.700 ;
        RECT 143.800 131.100 144.200 133.400 ;
        RECT 145.600 133.100 145.900 133.800 ;
        RECT 148.000 133.700 148.300 134.500 ;
        RECT 148.800 134.200 149.100 135.800 ;
        RECT 151.800 135.700 152.200 139.900 ;
        RECT 154.000 138.200 154.400 139.900 ;
        RECT 153.400 137.900 154.400 138.200 ;
        RECT 156.200 137.900 156.600 139.900 ;
        RECT 158.300 137.900 158.900 139.900 ;
        RECT 153.400 137.500 153.800 137.900 ;
        RECT 156.200 137.600 156.500 137.900 ;
        RECT 155.100 137.300 156.900 137.600 ;
        RECT 158.200 137.500 158.600 137.900 ;
        RECT 155.100 137.200 155.500 137.300 ;
        RECT 156.500 137.200 156.900 137.300 ;
        RECT 153.400 136.500 153.800 136.600 ;
        RECT 155.700 136.500 156.100 136.600 ;
        RECT 153.400 136.200 156.100 136.500 ;
        RECT 156.400 136.500 157.500 136.800 ;
        RECT 156.400 135.900 156.700 136.500 ;
        RECT 157.100 136.400 157.500 136.500 ;
        RECT 158.300 136.600 159.000 137.000 ;
        RECT 158.300 136.100 158.600 136.600 ;
        RECT 154.300 135.700 156.700 135.900 ;
        RECT 151.800 135.600 156.700 135.700 ;
        RECT 157.400 135.800 158.600 136.100 ;
        RECT 151.800 135.500 154.700 135.600 ;
        RECT 151.800 135.400 154.600 135.500 ;
        RECT 155.000 135.100 155.400 135.200 ;
        RECT 156.600 135.100 157.000 135.200 ;
        RECT 152.900 134.800 157.000 135.100 ;
        RECT 152.900 134.700 153.300 134.800 ;
        RECT 153.700 134.200 154.100 134.300 ;
        RECT 157.400 134.200 157.700 135.800 ;
        RECT 160.600 135.600 161.000 139.900 ;
        RECT 161.700 139.200 162.100 139.900 ;
        RECT 161.400 138.800 162.100 139.200 ;
        RECT 161.700 136.300 162.100 138.800 ;
        RECT 161.700 135.900 162.600 136.300 ;
        RECT 158.900 135.300 161.000 135.600 ;
        RECT 158.900 135.200 159.300 135.300 ;
        RECT 159.700 134.900 160.100 135.000 ;
        RECT 158.200 134.600 160.100 134.900 ;
        RECT 158.200 134.500 158.600 134.600 ;
        RECT 148.600 133.800 149.100 134.200 ;
        RECT 152.200 133.900 157.700 134.200 ;
        RECT 152.200 133.800 153.000 133.900 ;
        RECT 145.400 132.800 145.900 133.100 ;
        RECT 147.000 133.400 148.300 133.700 ;
        RECT 145.400 131.100 145.800 132.800 ;
        RECT 147.000 131.100 147.400 133.400 ;
        RECT 148.800 133.100 149.100 133.800 ;
        RECT 148.600 132.800 149.100 133.100 ;
        RECT 148.600 131.100 149.000 132.800 ;
        RECT 151.800 131.100 152.200 133.500 ;
        RECT 154.300 132.800 154.600 133.900 ;
        RECT 157.100 133.800 157.500 133.900 ;
        RECT 160.600 133.600 161.000 135.300 ;
        RECT 161.400 134.800 161.800 135.600 ;
        RECT 159.100 133.300 161.000 133.600 ;
        RECT 159.100 133.200 159.500 133.300 ;
        RECT 160.600 133.100 161.000 133.300 ;
        RECT 162.200 134.200 162.500 135.900 ;
        RECT 163.800 135.100 164.200 135.200 ;
        RECT 164.600 135.100 165.000 139.900 ;
        RECT 165.400 137.500 165.800 139.500 ;
        RECT 165.400 135.800 165.700 137.500 ;
        RECT 167.500 136.400 167.900 139.900 ;
        RECT 167.500 136.100 168.300 136.400 ;
        RECT 165.400 135.500 167.300 135.800 ;
        RECT 163.800 134.800 165.000 135.100 ;
        RECT 162.200 133.800 162.600 134.200 ;
        RECT 161.400 133.100 161.800 133.200 ;
        RECT 160.600 132.800 161.800 133.100 ;
        RECT 153.400 132.100 153.800 132.500 ;
        RECT 154.200 132.400 154.600 132.800 ;
        RECT 155.100 132.700 155.500 132.800 ;
        RECT 155.100 132.400 156.500 132.700 ;
        RECT 156.200 132.100 156.500 132.400 ;
        RECT 158.200 132.100 158.600 132.500 ;
        RECT 153.400 131.800 154.400 132.100 ;
        RECT 154.000 131.100 154.400 131.800 ;
        RECT 156.200 131.100 156.600 132.100 ;
        RECT 158.200 131.800 158.900 132.100 ;
        RECT 158.300 131.100 158.900 131.800 ;
        RECT 160.600 131.100 161.000 132.800 ;
        RECT 162.200 132.100 162.500 133.800 ;
        RECT 163.000 132.400 163.400 133.200 ;
        RECT 163.800 132.400 164.200 133.200 ;
        RECT 162.200 131.100 162.600 132.100 ;
        RECT 164.600 131.100 165.000 134.800 ;
        RECT 165.400 134.400 165.800 135.200 ;
        RECT 166.200 134.400 166.600 135.200 ;
        RECT 167.000 134.500 167.300 135.500 ;
        RECT 167.000 134.100 167.700 134.500 ;
        RECT 168.000 134.200 168.300 136.100 ;
        RECT 170.200 135.800 170.600 136.600 ;
        RECT 168.600 134.800 169.000 135.600 ;
        RECT 167.000 133.900 167.500 134.100 ;
        RECT 165.400 133.600 167.500 133.900 ;
        RECT 168.000 133.800 169.000 134.200 ;
        RECT 165.400 132.500 165.700 133.600 ;
        RECT 168.000 133.500 168.300 133.800 ;
        RECT 167.900 133.300 168.300 133.500 ;
        RECT 167.500 133.000 168.300 133.300 ;
        RECT 171.000 133.100 171.400 139.900 ;
        RECT 173.000 136.800 173.400 137.200 ;
        RECT 173.000 136.200 173.300 136.800 ;
        RECT 173.700 136.200 174.100 139.900 ;
        RECT 175.800 137.900 176.200 139.900 ;
        RECT 175.900 137.800 176.200 137.900 ;
        RECT 177.400 137.900 177.800 139.900 ;
        RECT 177.400 137.800 177.700 137.900 ;
        RECT 175.900 137.500 177.700 137.800 ;
        RECT 175.900 136.200 176.200 137.500 ;
        RECT 176.600 136.400 177.000 137.200 ;
        RECT 172.600 135.900 173.300 136.200 ;
        RECT 173.600 135.900 174.100 136.200 ;
        RECT 172.600 135.800 173.000 135.900 ;
        RECT 171.800 135.100 172.200 135.200 ;
        RECT 173.600 135.100 173.900 135.900 ;
        RECT 175.800 135.800 176.200 136.200 ;
        RECT 171.800 134.800 173.900 135.100 ;
        RECT 173.600 134.200 173.900 134.800 ;
        RECT 174.200 134.400 174.600 135.200 ;
        RECT 175.900 134.200 176.200 135.800 ;
        RECT 178.200 135.400 178.600 136.200 ;
        RECT 177.000 134.800 177.800 135.200 ;
        RECT 179.000 135.100 179.400 135.200 ;
        RECT 179.800 135.100 180.200 139.900 ;
        RECT 179.000 134.800 180.200 135.100 ;
        RECT 180.600 136.100 181.000 136.600 ;
        RECT 181.400 136.100 181.800 139.900 ;
        RECT 180.600 135.900 181.800 136.100 ;
        RECT 183.000 137.900 183.400 139.900 ;
        RECT 180.600 135.800 181.700 135.900 ;
        RECT 183.000 135.800 183.300 137.900 ;
        RECT 185.000 136.800 185.400 137.200 ;
        RECT 185.000 136.200 185.300 136.800 ;
        RECT 185.700 136.200 186.100 139.900 ;
        RECT 184.600 135.900 185.300 136.200 ;
        RECT 185.600 135.900 186.100 136.200 ;
        RECT 184.600 135.800 185.000 135.900 ;
        RECT 180.600 135.200 180.900 135.800 ;
        RECT 181.400 135.200 181.700 135.800 ;
        RECT 182.100 135.500 183.300 135.800 ;
        RECT 180.600 134.800 181.000 135.200 ;
        RECT 181.400 134.800 181.800 135.200 ;
        RECT 172.600 133.800 173.900 134.200 ;
        RECT 175.000 134.100 175.400 134.200 ;
        RECT 174.600 133.800 175.400 134.100 ;
        RECT 175.900 134.100 176.700 134.200 ;
        RECT 175.900 133.900 176.800 134.100 ;
        RECT 172.700 133.100 173.000 133.800 ;
        RECT 174.600 133.600 175.000 133.800 ;
        RECT 173.500 133.100 175.300 133.300 ;
        RECT 165.400 131.500 165.800 132.500 ;
        RECT 167.500 132.200 167.900 133.000 ;
        RECT 170.500 132.800 171.400 133.100 ;
        RECT 170.500 132.200 170.900 132.800 ;
        RECT 167.500 131.800 168.200 132.200 ;
        RECT 170.200 131.800 170.900 132.200 ;
        RECT 167.500 131.500 167.900 131.800 ;
        RECT 170.500 131.100 170.900 131.800 ;
        RECT 172.600 131.100 173.000 133.100 ;
        RECT 173.400 133.000 175.400 133.100 ;
        RECT 173.400 131.100 173.800 133.000 ;
        RECT 175.000 131.100 175.400 133.000 ;
        RECT 176.400 131.100 176.800 133.900 ;
        RECT 179.000 133.400 179.400 134.200 ;
        RECT 179.800 134.100 180.200 134.800 ;
        RECT 180.600 134.100 181.000 134.200 ;
        RECT 179.800 133.800 181.000 134.100 ;
        RECT 179.800 133.100 180.200 133.800 ;
        RECT 181.400 133.100 181.700 134.800 ;
        RECT 182.100 133.800 182.400 135.500 ;
        RECT 185.600 135.200 185.900 135.900 ;
        RECT 187.800 135.800 188.200 136.600 ;
        RECT 183.000 134.800 183.400 135.200 ;
        RECT 185.400 134.800 185.900 135.200 ;
        RECT 183.000 134.400 183.300 134.800 ;
        RECT 182.800 134.100 183.300 134.400 ;
        RECT 182.800 134.000 183.200 134.100 ;
        RECT 183.800 133.800 184.200 134.600 ;
        RECT 185.600 134.200 185.900 134.800 ;
        RECT 186.200 134.400 186.600 135.200 ;
        RECT 184.600 133.800 185.900 134.200 ;
        RECT 187.000 134.100 187.400 134.200 ;
        RECT 188.600 134.100 189.000 139.900 ;
        RECT 190.200 135.800 190.600 136.600 ;
        RECT 186.600 133.800 189.000 134.100 ;
        RECT 182.000 133.700 182.400 133.800 ;
        RECT 182.000 133.500 183.500 133.700 ;
        RECT 182.000 133.400 184.100 133.500 ;
        RECT 183.200 133.200 184.100 133.400 ;
        RECT 183.800 133.100 184.100 133.200 ;
        RECT 184.700 133.100 185.000 133.800 ;
        RECT 186.600 133.600 187.000 133.800 ;
        RECT 185.500 133.100 187.300 133.300 ;
        RECT 188.600 133.100 189.000 133.800 ;
        RECT 189.400 133.400 189.800 134.200 ;
        RECT 191.000 133.100 191.400 139.900 ;
        RECT 192.600 137.900 193.000 139.900 ;
        RECT 192.700 137.800 193.000 137.900 ;
        RECT 194.200 137.900 194.600 139.900 ;
        RECT 194.200 137.800 194.500 137.900 ;
        RECT 192.700 137.500 194.500 137.800 ;
        RECT 192.700 136.200 193.000 137.500 ;
        RECT 193.400 136.400 193.800 137.200 ;
        RECT 192.600 135.800 193.000 136.200 ;
        RECT 192.700 134.200 193.000 135.800 ;
        RECT 195.000 135.400 195.400 136.200 ;
        RECT 195.800 135.900 196.200 139.900 ;
        RECT 196.600 136.200 197.000 139.900 ;
        RECT 198.200 136.200 198.600 139.900 ;
        RECT 196.600 135.900 198.600 136.200 ;
        RECT 199.000 136.200 199.400 139.900 ;
        RECT 199.800 136.200 200.200 136.300 ;
        RECT 201.200 136.200 202.000 139.900 ;
        RECT 199.000 135.900 200.200 136.200 ;
        RECT 201.000 135.900 202.000 136.200 ;
        RECT 203.100 136.200 203.500 136.300 ;
        RECT 203.800 136.200 204.200 139.900 ;
        RECT 203.100 135.900 204.200 136.200 ;
        RECT 195.900 135.200 196.200 135.900 ;
        RECT 201.000 135.200 201.300 135.900 ;
        RECT 203.100 135.600 203.400 135.900 ;
        RECT 201.700 135.300 203.400 135.600 ;
        RECT 201.700 135.200 202.100 135.300 ;
        RECT 193.800 134.800 194.600 135.200 ;
        RECT 195.800 134.900 197.000 135.200 ;
        RECT 195.800 134.800 196.200 134.900 ;
        RECT 191.800 133.400 192.200 134.200 ;
        RECT 192.700 134.100 193.500 134.200 ;
        RECT 195.800 134.100 196.200 134.200 ;
        RECT 196.700 134.100 197.000 134.900 ;
        RECT 200.600 134.900 201.300 135.200 ;
        RECT 202.800 134.900 203.200 135.000 ;
        RECT 200.600 134.800 201.500 134.900 ;
        RECT 201.000 134.600 201.500 134.800 ;
        RECT 192.700 133.900 193.600 134.100 ;
        RECT 179.800 132.800 180.700 133.100 ;
        RECT 180.300 131.100 180.700 132.800 ;
        RECT 181.400 132.600 182.100 133.100 ;
        RECT 181.700 131.100 182.100 132.600 ;
        RECT 183.800 131.100 184.200 133.100 ;
        RECT 184.600 131.100 185.000 133.100 ;
        RECT 185.400 133.000 187.400 133.100 ;
        RECT 185.400 131.100 185.800 133.000 ;
        RECT 187.000 131.100 187.400 133.000 ;
        RECT 188.100 132.800 189.000 133.100 ;
        RECT 190.500 132.800 191.400 133.100 ;
        RECT 188.100 131.100 188.500 132.800 ;
        RECT 190.500 131.100 190.900 132.800 ;
        RECT 193.200 131.100 193.600 133.900 ;
        RECT 195.800 133.800 197.000 134.100 ;
        RECT 197.400 133.800 197.800 134.600 ;
        RECT 199.000 133.800 199.800 134.200 ;
        RECT 200.400 133.800 200.800 134.200 ;
        RECT 195.800 132.800 196.200 133.200 ;
        RECT 196.700 133.100 197.000 133.800 ;
        RECT 200.500 133.600 200.800 133.800 ;
        RECT 199.800 133.400 200.200 133.500 ;
        RECT 195.900 132.400 196.300 132.800 ;
        RECT 196.600 131.100 197.000 133.100 ;
        RECT 199.000 133.100 200.200 133.400 ;
        RECT 200.500 133.200 200.900 133.600 ;
        RECT 199.000 131.100 199.400 133.100 ;
        RECT 201.200 132.900 201.500 134.600 ;
        RECT 201.900 134.600 203.200 134.900 ;
        RECT 201.900 134.300 202.200 134.600 ;
        RECT 201.800 133.900 202.200 134.300 ;
        RECT 203.400 134.100 204.200 134.200 ;
        RECT 204.600 134.100 205.000 134.200 ;
        RECT 202.500 133.800 205.000 134.100 ;
        RECT 202.500 133.600 202.800 133.800 ;
        RECT 201.800 133.300 202.800 133.600 ;
        RECT 203.100 133.400 203.500 133.500 ;
        RECT 201.800 133.200 202.600 133.300 ;
        RECT 203.100 133.100 204.200 133.400 ;
        RECT 201.200 131.100 202.000 132.900 ;
        RECT 203.800 131.100 204.200 133.100 ;
        RECT 0.600 127.500 1.000 129.900 ;
        RECT 2.800 129.200 3.200 129.900 ;
        RECT 2.200 128.900 3.200 129.200 ;
        RECT 5.000 128.900 5.400 129.900 ;
        RECT 7.100 129.200 7.700 129.900 ;
        RECT 7.000 128.900 7.700 129.200 ;
        RECT 2.200 128.500 2.600 128.900 ;
        RECT 5.000 128.600 5.300 128.900 ;
        RECT 3.000 127.800 3.400 128.600 ;
        RECT 3.900 128.300 5.300 128.600 ;
        RECT 7.000 128.500 7.400 128.900 ;
        RECT 3.900 128.200 4.300 128.300 ;
        RECT 9.400 128.100 9.800 129.900 ;
        RECT 10.200 128.100 10.600 128.600 ;
        RECT 9.400 127.800 10.600 128.100 ;
        RECT 1.000 127.100 1.800 127.200 ;
        RECT 3.100 127.100 3.400 127.800 ;
        RECT 7.900 127.700 8.300 127.800 ;
        RECT 9.400 127.700 9.800 127.800 ;
        RECT 7.900 127.400 9.800 127.700 ;
        RECT 5.900 127.100 6.300 127.200 ;
        RECT 1.000 126.800 6.500 127.100 ;
        RECT 2.500 126.700 2.900 126.800 ;
        RECT 1.700 126.200 2.100 126.300 ;
        RECT 1.700 126.100 4.200 126.200 ;
        RECT 5.400 126.100 5.800 126.200 ;
        RECT 1.700 125.900 5.800 126.100 ;
        RECT 3.800 125.800 5.800 125.900 ;
        RECT 0.600 125.500 3.400 125.600 ;
        RECT 0.600 125.400 3.500 125.500 ;
        RECT 0.600 125.300 5.500 125.400 ;
        RECT 0.600 121.100 1.000 125.300 ;
        RECT 3.100 125.100 5.500 125.300 ;
        RECT 2.200 124.500 4.900 124.800 ;
        RECT 2.200 124.400 2.600 124.500 ;
        RECT 4.500 124.400 4.900 124.500 ;
        RECT 5.200 124.500 5.500 125.100 ;
        RECT 6.200 125.200 6.500 126.800 ;
        RECT 7.000 126.400 7.400 126.500 ;
        RECT 7.000 126.100 8.900 126.400 ;
        RECT 8.500 126.000 8.900 126.100 ;
        RECT 7.700 125.700 8.100 125.800 ;
        RECT 9.400 125.700 9.800 127.400 ;
        RECT 7.700 125.400 9.800 125.700 ;
        RECT 6.200 124.900 7.400 125.200 ;
        RECT 5.900 124.500 6.300 124.600 ;
        RECT 5.200 124.200 6.300 124.500 ;
        RECT 7.100 124.400 7.400 124.900 ;
        RECT 7.100 124.000 7.800 124.400 ;
        RECT 3.900 123.700 4.300 123.800 ;
        RECT 5.300 123.700 5.700 123.800 ;
        RECT 2.200 123.100 2.600 123.500 ;
        RECT 3.900 123.400 5.700 123.700 ;
        RECT 5.000 123.100 5.300 123.400 ;
        RECT 7.000 123.100 7.400 123.500 ;
        RECT 2.200 122.800 3.200 123.100 ;
        RECT 2.800 121.100 3.200 122.800 ;
        RECT 5.000 121.100 5.400 123.100 ;
        RECT 7.100 121.100 7.700 123.100 ;
        RECT 9.400 121.100 9.800 125.400 ;
        RECT 11.000 121.100 11.400 129.900 ;
        RECT 13.700 128.000 14.100 129.500 ;
        RECT 15.800 128.500 16.200 129.500 ;
        RECT 13.300 127.700 14.100 128.000 ;
        RECT 13.300 127.500 13.700 127.700 ;
        RECT 13.300 127.200 13.600 127.500 ;
        RECT 15.900 127.400 16.200 128.500 ;
        RECT 16.600 127.500 17.000 129.900 ;
        RECT 18.800 129.200 19.200 129.900 ;
        RECT 18.200 128.900 19.200 129.200 ;
        RECT 21.000 128.900 21.400 129.900 ;
        RECT 23.100 129.200 23.700 129.900 ;
        RECT 23.000 128.900 23.700 129.200 ;
        RECT 18.200 128.500 18.600 128.900 ;
        RECT 21.000 128.600 21.300 128.900 ;
        RECT 19.000 128.200 19.400 128.600 ;
        RECT 19.900 128.300 21.300 128.600 ;
        RECT 23.000 128.500 23.400 128.900 ;
        RECT 19.900 128.200 20.300 128.300 ;
        RECT 12.600 126.800 13.600 127.200 ;
        RECT 14.100 127.100 16.200 127.400 ;
        RECT 17.000 127.100 17.800 127.200 ;
        RECT 19.100 127.100 19.400 128.200 ;
        RECT 23.900 127.700 24.300 127.800 ;
        RECT 25.400 127.700 25.800 129.900 ;
        RECT 26.200 128.000 26.600 129.900 ;
        RECT 27.800 128.000 28.200 129.900 ;
        RECT 26.200 127.900 28.200 128.000 ;
        RECT 28.600 127.900 29.000 129.900 ;
        RECT 29.700 128.200 30.100 129.900 ;
        RECT 29.700 127.900 30.600 128.200 ;
        RECT 26.300 127.700 28.100 127.900 ;
        RECT 23.900 127.400 25.800 127.700 ;
        RECT 21.900 127.100 22.300 127.200 ;
        RECT 14.100 126.900 14.600 127.100 ;
        RECT 12.600 125.400 13.000 126.200 ;
        RECT 13.300 124.900 13.600 126.800 ;
        RECT 13.900 126.500 14.600 126.900 ;
        RECT 17.000 126.800 22.500 127.100 ;
        RECT 18.500 126.700 18.900 126.800 ;
        RECT 14.300 125.500 14.600 126.500 ;
        RECT 15.000 125.800 15.400 126.600 ;
        RECT 15.800 125.800 16.200 126.600 ;
        RECT 17.700 126.200 18.100 126.300 ;
        RECT 17.700 125.900 20.200 126.200 ;
        RECT 19.800 125.800 20.200 125.900 ;
        RECT 16.600 125.500 19.400 125.600 ;
        RECT 14.300 125.200 16.200 125.500 ;
        RECT 13.300 124.600 14.100 124.900 ;
        RECT 13.700 121.100 14.100 124.600 ;
        RECT 15.900 123.500 16.200 125.200 ;
        RECT 15.800 121.500 16.200 123.500 ;
        RECT 16.600 125.400 19.500 125.500 ;
        RECT 16.600 125.300 21.500 125.400 ;
        RECT 16.600 121.100 17.000 125.300 ;
        RECT 19.100 125.100 21.500 125.300 ;
        RECT 18.200 124.500 20.900 124.800 ;
        RECT 18.200 124.400 18.600 124.500 ;
        RECT 20.500 124.400 20.900 124.500 ;
        RECT 21.200 124.500 21.500 125.100 ;
        RECT 22.200 125.200 22.500 126.800 ;
        RECT 23.000 126.400 23.400 126.500 ;
        RECT 23.000 126.100 24.900 126.400 ;
        RECT 24.500 126.000 24.900 126.100 ;
        RECT 23.700 125.700 24.100 125.800 ;
        RECT 25.400 125.700 25.800 127.400 ;
        RECT 26.600 127.200 27.000 127.400 ;
        RECT 28.600 127.200 28.900 127.900 ;
        RECT 26.200 126.900 27.000 127.200 ;
        RECT 26.200 126.800 26.600 126.900 ;
        RECT 27.700 126.800 29.000 127.200 ;
        RECT 27.000 125.800 27.400 126.600 ;
        RECT 23.700 125.400 25.800 125.700 ;
        RECT 22.200 124.900 23.400 125.200 ;
        RECT 21.900 124.500 22.300 124.600 ;
        RECT 21.200 124.200 22.300 124.500 ;
        RECT 23.100 124.400 23.400 124.900 ;
        RECT 23.100 124.000 23.800 124.400 ;
        RECT 19.900 123.700 20.300 123.800 ;
        RECT 21.300 123.700 21.700 123.800 ;
        RECT 18.200 123.100 18.600 123.500 ;
        RECT 19.900 123.400 21.700 123.700 ;
        RECT 21.000 123.100 21.300 123.400 ;
        RECT 23.000 123.100 23.400 123.500 ;
        RECT 18.200 122.800 19.200 123.100 ;
        RECT 18.800 121.100 19.200 122.800 ;
        RECT 21.000 121.100 21.400 123.100 ;
        RECT 23.100 121.100 23.700 123.100 ;
        RECT 25.400 121.100 25.800 125.400 ;
        RECT 27.700 125.200 28.000 126.800 ;
        RECT 30.200 126.100 30.600 127.900 ;
        RECT 27.000 124.800 28.000 125.200 ;
        RECT 28.600 125.800 30.600 126.100 ;
        RECT 31.000 126.800 31.400 127.600 ;
        RECT 31.800 127.500 32.200 129.900 ;
        RECT 34.000 129.200 34.400 129.900 ;
        RECT 33.400 128.900 34.400 129.200 ;
        RECT 36.200 128.900 36.600 129.900 ;
        RECT 38.300 129.200 38.900 129.900 ;
        RECT 38.200 128.900 38.900 129.200 ;
        RECT 33.400 128.500 33.800 128.900 ;
        RECT 36.200 128.600 36.500 128.900 ;
        RECT 34.200 128.200 34.600 128.600 ;
        RECT 35.100 128.300 36.500 128.600 ;
        RECT 38.200 128.500 38.600 128.900 ;
        RECT 35.100 128.200 35.500 128.300 ;
        RECT 32.200 127.100 33.000 127.200 ;
        RECT 34.300 127.100 34.600 128.200 ;
        RECT 39.100 127.700 39.500 127.800 ;
        RECT 40.600 127.700 41.000 129.900 ;
        RECT 42.700 129.200 43.100 129.900 ;
        RECT 42.200 128.800 43.100 129.200 ;
        RECT 42.700 128.200 43.100 128.800 ;
        RECT 39.100 127.400 41.000 127.700 ;
        RECT 42.200 127.900 43.100 128.200 ;
        RECT 43.800 128.000 44.200 129.900 ;
        RECT 45.400 128.000 45.800 129.900 ;
        RECT 43.800 127.900 45.800 128.000 ;
        RECT 46.200 127.900 46.600 129.900 ;
        RECT 47.000 128.000 47.400 129.900 ;
        RECT 48.600 129.600 50.600 129.900 ;
        RECT 48.600 128.000 49.000 129.600 ;
        RECT 47.000 127.900 49.000 128.000 ;
        RECT 49.400 127.900 49.800 129.300 ;
        RECT 50.200 127.900 50.600 129.600 ;
        RECT 54.200 127.900 54.600 129.900 ;
        RECT 54.900 128.200 55.300 128.600 ;
        RECT 37.100 127.100 37.500 127.200 ;
        RECT 32.200 126.800 37.700 127.100 ;
        RECT 31.000 126.200 31.300 126.800 ;
        RECT 33.700 126.700 34.100 126.800 ;
        RECT 32.900 126.200 33.300 126.300 ;
        RECT 37.400 126.200 37.700 126.800 ;
        RECT 38.200 126.400 38.600 126.500 ;
        RECT 31.000 125.800 31.400 126.200 ;
        RECT 32.900 126.100 35.400 126.200 ;
        RECT 35.800 126.100 36.200 126.200 ;
        RECT 32.900 125.900 36.200 126.100 ;
        RECT 35.000 125.800 36.200 125.900 ;
        RECT 37.400 125.800 37.800 126.200 ;
        RECT 38.200 126.100 40.100 126.400 ;
        RECT 39.700 126.000 40.100 126.100 ;
        RECT 28.600 125.200 28.900 125.800 ;
        RECT 28.600 125.100 29.000 125.200 ;
        RECT 28.300 124.800 29.000 125.100 ;
        RECT 27.500 121.100 27.900 124.800 ;
        RECT 28.300 124.200 28.600 124.800 ;
        RECT 29.400 124.400 29.800 125.200 ;
        RECT 28.200 123.800 28.600 124.200 ;
        RECT 30.200 121.100 30.600 125.800 ;
        RECT 31.800 125.500 34.600 125.600 ;
        RECT 31.800 125.400 34.700 125.500 ;
        RECT 31.800 125.300 36.700 125.400 ;
        RECT 31.800 121.100 32.200 125.300 ;
        RECT 34.300 125.100 36.700 125.300 ;
        RECT 33.400 124.500 36.100 124.800 ;
        RECT 33.400 124.400 33.800 124.500 ;
        RECT 35.700 124.400 36.100 124.500 ;
        RECT 36.400 124.500 36.700 125.100 ;
        RECT 37.400 125.200 37.700 125.800 ;
        RECT 38.900 125.700 39.300 125.800 ;
        RECT 40.600 125.700 41.000 127.400 ;
        RECT 41.400 126.800 41.800 127.600 ;
        RECT 38.900 125.400 41.000 125.700 ;
        RECT 37.400 124.900 38.600 125.200 ;
        RECT 37.100 124.500 37.500 124.600 ;
        RECT 36.400 124.200 37.500 124.500 ;
        RECT 38.300 124.400 38.600 124.900 ;
        RECT 38.300 124.000 39.000 124.400 ;
        RECT 40.600 124.100 41.000 125.400 ;
        RECT 41.400 124.100 41.800 124.200 ;
        RECT 40.600 123.800 41.800 124.100 ;
        RECT 35.100 123.700 35.500 123.800 ;
        RECT 36.500 123.700 36.900 123.800 ;
        RECT 33.400 123.100 33.800 123.500 ;
        RECT 35.100 123.400 36.900 123.700 ;
        RECT 36.200 123.100 36.500 123.400 ;
        RECT 38.200 123.100 38.600 123.500 ;
        RECT 33.400 122.800 34.400 123.100 ;
        RECT 34.000 121.100 34.400 122.800 ;
        RECT 36.200 121.100 36.600 123.100 ;
        RECT 38.300 121.100 38.900 123.100 ;
        RECT 40.600 121.100 41.000 123.800 ;
        RECT 42.200 121.100 42.600 127.900 ;
        RECT 43.900 127.700 45.700 127.900 ;
        RECT 44.200 127.200 44.600 127.400 ;
        RECT 46.200 127.200 46.500 127.900 ;
        RECT 47.100 127.700 48.900 127.900 ;
        RECT 47.400 127.200 47.800 127.400 ;
        RECT 49.500 127.200 49.800 127.900 ;
        RECT 43.800 126.900 44.600 127.200 ;
        RECT 43.800 126.800 44.200 126.900 ;
        RECT 45.300 126.800 46.600 127.200 ;
        RECT 47.000 126.900 47.800 127.200 ;
        RECT 48.600 126.900 49.800 127.200 ;
        RECT 47.000 126.800 47.400 126.900 ;
        RECT 48.600 126.800 49.000 126.900 ;
        RECT 44.600 125.800 45.000 126.600 ;
        RECT 43.000 124.400 43.400 125.200 ;
        RECT 45.300 125.100 45.600 126.800 ;
        RECT 47.800 125.800 48.200 126.600 ;
        RECT 46.200 125.100 46.600 125.200 ;
        RECT 48.600 125.100 48.900 126.800 ;
        RECT 49.400 125.800 49.800 126.600 ;
        RECT 50.200 126.400 50.600 127.200 ;
        RECT 53.400 126.400 53.800 127.200 ;
        RECT 51.800 126.100 52.200 126.200 ;
        RECT 52.600 126.100 53.000 126.200 ;
        RECT 54.200 126.100 54.500 127.900 ;
        RECT 55.000 127.800 55.400 128.200 ;
        RECT 55.800 127.900 56.200 129.900 ;
        RECT 56.600 128.000 57.000 129.900 ;
        RECT 58.200 128.000 58.600 129.900 ;
        RECT 59.300 128.200 59.700 129.900 ;
        RECT 56.600 127.900 58.600 128.000 ;
        RECT 55.900 127.200 56.200 127.900 ;
        RECT 56.700 127.700 58.500 127.900 ;
        RECT 59.000 127.800 60.200 128.200 ;
        RECT 61.400 127.800 61.800 128.600 ;
        RECT 57.800 127.200 58.200 127.400 ;
        RECT 55.800 126.800 57.100 127.200 ;
        RECT 57.800 126.900 58.600 127.200 ;
        RECT 58.200 126.800 58.600 126.900 ;
        RECT 55.000 126.100 55.400 126.200 ;
        RECT 51.800 125.800 53.400 126.100 ;
        RECT 54.200 125.800 55.400 126.100 ;
        RECT 53.000 125.600 53.400 125.800 ;
        RECT 55.000 125.100 55.300 125.800 ;
        RECT 56.800 125.200 57.100 126.800 ;
        RECT 57.400 125.800 57.800 126.600 ;
        RECT 55.800 125.100 56.200 125.200 ;
        RECT 45.100 124.800 45.600 125.100 ;
        RECT 45.900 124.800 46.600 125.100 ;
        RECT 45.100 121.100 45.500 124.800 ;
        RECT 45.900 124.200 46.200 124.800 ;
        RECT 45.800 123.800 46.200 124.200 ;
        RECT 48.300 121.100 49.300 125.100 ;
        RECT 52.600 124.800 54.600 125.100 ;
        RECT 52.600 121.100 53.000 124.800 ;
        RECT 54.200 121.100 54.600 124.800 ;
        RECT 55.000 121.100 55.400 125.100 ;
        RECT 55.800 124.800 56.500 125.100 ;
        RECT 56.800 124.800 57.800 125.200 ;
        RECT 56.200 124.200 56.500 124.800 ;
        RECT 56.200 123.800 56.600 124.200 ;
        RECT 56.900 121.100 57.300 124.800 ;
        RECT 59.000 124.400 59.400 125.200 ;
        RECT 59.800 121.100 60.200 127.800 ;
        RECT 60.600 126.800 61.000 127.600 ;
        RECT 62.200 121.100 62.600 129.900 ;
        RECT 63.000 127.900 63.400 129.900 ;
        RECT 63.800 128.000 64.200 129.900 ;
        RECT 65.400 128.000 65.800 129.900 ;
        RECT 63.800 127.900 65.800 128.000 ;
        RECT 66.200 128.000 66.600 129.900 ;
        RECT 67.800 128.000 68.200 129.900 ;
        RECT 66.200 127.900 68.200 128.000 ;
        RECT 68.600 127.900 69.000 129.900 ;
        RECT 69.400 128.000 69.800 129.900 ;
        RECT 71.000 128.000 71.400 129.900 ;
        RECT 69.400 127.900 71.400 128.000 ;
        RECT 71.800 127.900 72.200 129.900 ;
        RECT 63.100 127.200 63.400 127.900 ;
        RECT 63.900 127.700 65.700 127.900 ;
        RECT 66.300 127.700 68.100 127.900 ;
        RECT 65.000 127.200 65.400 127.400 ;
        RECT 66.600 127.200 67.000 127.400 ;
        RECT 68.600 127.200 68.900 127.900 ;
        RECT 69.500 127.700 71.300 127.900 ;
        RECT 69.800 127.200 70.200 127.400 ;
        RECT 71.800 127.200 72.100 127.900 ;
        RECT 72.600 127.700 73.000 129.900 ;
        RECT 74.700 129.200 75.300 129.900 ;
        RECT 74.700 128.900 75.400 129.200 ;
        RECT 77.000 128.900 77.400 129.900 ;
        RECT 79.200 129.200 79.600 129.900 ;
        RECT 79.200 128.900 80.200 129.200 ;
        RECT 75.000 128.500 75.400 128.900 ;
        RECT 77.100 128.600 77.400 128.900 ;
        RECT 77.100 128.300 78.500 128.600 ;
        RECT 78.100 128.200 78.500 128.300 ;
        RECT 79.000 128.200 79.400 128.600 ;
        RECT 79.800 128.500 80.200 128.900 ;
        RECT 74.100 127.700 74.500 127.800 ;
        RECT 72.600 127.400 74.500 127.700 ;
        RECT 63.000 126.800 64.300 127.200 ;
        RECT 65.000 126.900 65.800 127.200 ;
        RECT 65.400 126.800 65.800 126.900 ;
        RECT 66.200 126.900 67.000 127.200 ;
        RECT 66.200 126.800 66.600 126.900 ;
        RECT 67.700 126.800 69.000 127.200 ;
        RECT 69.400 126.900 70.200 127.200 ;
        RECT 69.400 126.800 69.800 126.900 ;
        RECT 70.900 126.800 72.200 127.200 ;
        RECT 64.000 126.200 64.300 126.800 ;
        RECT 63.800 125.800 64.300 126.200 ;
        RECT 64.600 125.800 65.000 126.600 ;
        RECT 67.000 125.800 67.400 126.600 ;
        RECT 63.000 125.100 63.400 125.200 ;
        RECT 64.000 125.100 64.300 125.800 ;
        RECT 67.700 125.100 68.000 126.800 ;
        RECT 70.200 125.800 70.600 126.600 ;
        RECT 70.900 126.200 71.200 126.800 ;
        RECT 70.900 125.800 71.400 126.200 ;
        RECT 68.600 125.100 69.000 125.200 ;
        RECT 70.900 125.100 71.200 125.800 ;
        RECT 72.600 125.700 73.000 127.400 ;
        RECT 76.100 127.100 76.500 127.200 ;
        RECT 78.200 127.100 78.600 127.200 ;
        RECT 79.000 127.100 79.300 128.200 ;
        RECT 81.400 127.500 81.800 129.900 ;
        RECT 82.200 127.900 82.600 129.900 ;
        RECT 83.000 128.000 83.400 129.900 ;
        RECT 84.600 128.000 85.000 129.900 ;
        RECT 83.000 127.900 85.000 128.000 ;
        RECT 86.200 128.900 86.600 129.900 ;
        RECT 82.300 127.200 82.600 127.900 ;
        RECT 83.100 127.700 84.900 127.900 ;
        RECT 84.200 127.200 84.600 127.400 ;
        RECT 86.200 127.200 86.500 128.900 ;
        RECT 87.000 127.800 87.400 128.600 ;
        RECT 80.600 127.100 81.400 127.200 ;
        RECT 75.900 126.800 81.400 127.100 ;
        RECT 82.200 126.800 83.500 127.200 ;
        RECT 84.200 126.900 85.000 127.200 ;
        RECT 84.600 126.800 85.000 126.900 ;
        RECT 86.200 126.800 86.600 127.200 ;
        RECT 75.000 126.400 75.400 126.500 ;
        RECT 73.500 126.100 75.400 126.400 ;
        RECT 73.500 126.000 73.900 126.100 ;
        RECT 74.300 125.700 74.700 125.800 ;
        RECT 72.600 125.400 74.700 125.700 ;
        RECT 71.800 125.100 72.200 125.200 ;
        RECT 63.000 124.800 63.700 125.100 ;
        RECT 64.000 124.800 64.500 125.100 ;
        RECT 63.400 124.200 63.700 124.800 ;
        RECT 63.400 123.800 63.800 124.200 ;
        RECT 64.100 121.100 64.500 124.800 ;
        RECT 67.500 124.800 68.000 125.100 ;
        RECT 68.300 124.800 69.000 125.100 ;
        RECT 70.700 124.800 71.200 125.100 ;
        RECT 71.500 124.800 72.200 125.100 ;
        RECT 67.500 121.100 67.900 124.800 ;
        RECT 68.300 124.200 68.600 124.800 ;
        RECT 68.200 123.800 68.600 124.200 ;
        RECT 70.700 121.100 71.100 124.800 ;
        RECT 71.500 124.200 71.800 124.800 ;
        RECT 71.400 123.800 71.800 124.200 ;
        RECT 72.600 121.100 73.000 125.400 ;
        RECT 75.900 125.200 76.200 126.800 ;
        RECT 79.500 126.700 79.900 126.800 ;
        RECT 80.300 126.200 80.700 126.300 ;
        RECT 77.400 126.100 77.800 126.200 ;
        RECT 78.200 126.100 80.700 126.200 ;
        RECT 77.400 125.900 80.700 126.100 ;
        RECT 77.400 125.800 78.600 125.900 ;
        RECT 79.000 125.500 81.800 125.600 ;
        RECT 78.900 125.400 81.800 125.500 ;
        RECT 75.000 124.900 76.200 125.200 ;
        RECT 76.900 125.300 81.800 125.400 ;
        RECT 76.900 125.100 79.300 125.300 ;
        RECT 75.000 124.400 75.300 124.900 ;
        RECT 74.600 124.000 75.300 124.400 ;
        RECT 76.100 124.500 76.500 124.600 ;
        RECT 76.900 124.500 77.200 125.100 ;
        RECT 76.100 124.200 77.200 124.500 ;
        RECT 77.500 124.500 80.200 124.800 ;
        RECT 77.500 124.400 77.900 124.500 ;
        RECT 79.800 124.400 80.200 124.500 ;
        RECT 76.700 123.700 77.100 123.800 ;
        RECT 78.100 123.700 78.500 123.800 ;
        RECT 75.000 123.100 75.400 123.500 ;
        RECT 76.700 123.400 78.500 123.700 ;
        RECT 77.100 123.100 77.400 123.400 ;
        RECT 79.800 123.100 80.200 123.500 ;
        RECT 74.700 121.100 75.300 123.100 ;
        RECT 77.000 121.100 77.400 123.100 ;
        RECT 79.200 122.800 80.200 123.100 ;
        RECT 79.200 121.100 79.600 122.800 ;
        RECT 81.400 121.100 81.800 125.300 ;
        RECT 82.200 125.100 82.600 125.200 ;
        RECT 83.200 125.100 83.500 126.800 ;
        RECT 83.800 125.800 84.200 126.600 ;
        RECT 85.400 125.400 85.800 126.200 ;
        RECT 86.200 125.100 86.500 126.800 ;
        RECT 82.200 124.800 82.900 125.100 ;
        RECT 83.200 124.800 83.700 125.100 ;
        RECT 82.600 124.200 82.900 124.800 ;
        RECT 82.600 123.800 83.000 124.200 ;
        RECT 83.300 122.200 83.700 124.800 ;
        RECT 85.700 124.700 86.600 125.100 ;
        RECT 85.700 122.200 86.100 124.700 ;
        RECT 83.300 121.800 84.200 122.200 ;
        RECT 85.700 121.800 86.600 122.200 ;
        RECT 83.300 121.100 83.700 121.800 ;
        RECT 85.700 121.100 86.100 121.800 ;
        RECT 87.800 121.100 88.200 129.900 ;
        RECT 88.600 128.100 89.000 128.600 ;
        RECT 89.400 128.100 89.800 129.900 ;
        RECT 91.500 129.200 92.100 129.900 ;
        RECT 91.500 128.900 92.200 129.200 ;
        RECT 93.800 128.900 94.200 129.900 ;
        RECT 96.000 129.200 96.400 129.900 ;
        RECT 96.000 128.900 97.000 129.200 ;
        RECT 91.800 128.500 92.200 128.900 ;
        RECT 93.900 128.600 94.200 128.900 ;
        RECT 93.900 128.300 95.300 128.600 ;
        RECT 94.900 128.200 95.300 128.300 ;
        RECT 95.800 128.200 96.200 128.600 ;
        RECT 96.600 128.500 97.000 128.900 ;
        RECT 88.600 127.800 89.800 128.100 ;
        RECT 89.400 127.700 89.800 127.800 ;
        RECT 90.900 127.700 91.300 127.800 ;
        RECT 89.400 127.400 91.300 127.700 ;
        RECT 89.400 125.700 89.800 127.400 ;
        RECT 92.900 127.100 93.300 127.200 ;
        RECT 95.800 127.100 96.100 128.200 ;
        RECT 98.200 127.500 98.600 129.900 ;
        RECT 100.300 128.200 100.700 129.900 ;
        RECT 99.800 127.900 100.700 128.200 ;
        RECT 103.000 127.900 103.400 129.900 ;
        RECT 103.800 128.000 104.200 129.900 ;
        RECT 105.400 128.000 105.800 129.900 ;
        RECT 103.800 127.900 105.800 128.000 ;
        RECT 106.200 127.900 106.600 129.900 ;
        RECT 107.000 128.000 107.400 129.900 ;
        RECT 108.600 128.000 109.000 129.900 ;
        RECT 107.000 127.900 109.000 128.000 ;
        RECT 109.400 129.600 111.400 129.900 ;
        RECT 109.400 127.900 109.800 129.600 ;
        RECT 97.400 127.100 98.200 127.200 ;
        RECT 92.700 126.800 98.200 127.100 ;
        RECT 99.000 126.800 99.400 127.600 ;
        RECT 91.800 126.400 92.200 126.500 ;
        RECT 90.300 126.100 92.200 126.400 ;
        RECT 92.700 126.200 93.000 126.800 ;
        RECT 96.300 126.700 96.700 126.800 ;
        RECT 97.100 126.200 97.500 126.300 ;
        RECT 90.300 126.000 90.700 126.100 ;
        RECT 92.600 125.800 93.000 126.200 ;
        RECT 95.000 125.900 97.500 126.200 ;
        RECT 99.800 126.100 100.200 127.900 ;
        RECT 103.100 127.200 103.400 127.900 ;
        RECT 103.900 127.700 105.700 127.900 ;
        RECT 105.000 127.200 105.400 127.400 ;
        RECT 106.300 127.200 106.600 127.900 ;
        RECT 107.100 127.700 108.900 127.900 ;
        RECT 110.200 127.800 110.600 129.300 ;
        RECT 111.000 128.000 111.400 129.600 ;
        RECT 112.600 128.000 113.000 129.900 ;
        RECT 111.000 127.900 113.000 128.000 ;
        RECT 114.200 128.900 114.600 129.900 ;
        RECT 116.600 128.900 117.000 129.900 ;
        RECT 108.200 127.200 108.600 127.400 ;
        RECT 110.200 127.200 110.500 127.800 ;
        RECT 111.100 127.700 112.900 127.900 ;
        RECT 112.200 127.200 112.600 127.400 ;
        RECT 114.200 127.200 114.500 128.900 ;
        RECT 115.000 127.800 115.400 128.600 ;
        RECT 115.800 127.800 116.200 128.600 ;
        RECT 116.700 127.200 117.000 128.900 ;
        RECT 100.600 127.100 101.000 127.200 ;
        RECT 103.000 127.100 104.300 127.200 ;
        RECT 100.600 126.800 104.300 127.100 ;
        RECT 105.000 126.900 105.800 127.200 ;
        RECT 105.400 126.800 105.800 126.900 ;
        RECT 106.200 126.800 107.500 127.200 ;
        RECT 108.200 126.900 109.000 127.200 ;
        RECT 108.600 126.800 109.000 126.900 ;
        RECT 95.000 125.800 95.400 125.900 ;
        RECT 99.800 125.800 103.300 126.100 ;
        RECT 91.100 125.700 91.500 125.800 ;
        RECT 89.400 125.400 91.500 125.700 ;
        RECT 89.400 121.100 89.800 125.400 ;
        RECT 92.700 125.200 93.000 125.800 ;
        RECT 95.800 125.500 98.600 125.600 ;
        RECT 95.700 125.400 98.600 125.500 ;
        RECT 91.800 124.900 93.000 125.200 ;
        RECT 93.700 125.300 98.600 125.400 ;
        RECT 93.700 125.100 96.100 125.300 ;
        RECT 91.800 124.400 92.100 124.900 ;
        RECT 91.400 124.000 92.100 124.400 ;
        RECT 92.900 124.500 93.300 124.600 ;
        RECT 93.700 124.500 94.000 125.100 ;
        RECT 92.900 124.200 94.000 124.500 ;
        RECT 94.300 124.500 97.000 124.800 ;
        RECT 94.300 124.400 94.700 124.500 ;
        RECT 96.600 124.400 97.000 124.500 ;
        RECT 93.500 123.700 93.900 123.800 ;
        RECT 94.900 123.700 95.300 123.800 ;
        RECT 91.800 123.100 92.200 123.500 ;
        RECT 93.500 123.400 95.300 123.700 ;
        RECT 93.900 123.100 94.200 123.400 ;
        RECT 96.600 123.100 97.000 123.500 ;
        RECT 91.500 121.100 92.100 123.100 ;
        RECT 93.800 121.100 94.200 123.100 ;
        RECT 96.000 122.800 97.000 123.100 ;
        RECT 96.000 121.100 96.400 122.800 ;
        RECT 98.200 121.100 98.600 125.300 ;
        RECT 99.800 121.100 100.200 125.800 ;
        RECT 103.000 125.200 103.300 125.800 ;
        RECT 100.600 124.400 101.000 125.200 ;
        RECT 103.000 125.100 103.400 125.200 ;
        RECT 104.000 125.100 104.300 126.800 ;
        RECT 104.600 125.800 105.000 126.600 ;
        RECT 106.200 125.100 106.600 125.200 ;
        RECT 107.200 125.100 107.500 126.800 ;
        RECT 107.800 125.800 108.200 126.600 ;
        RECT 109.400 126.400 109.800 127.200 ;
        RECT 110.200 126.900 111.400 127.200 ;
        RECT 112.200 127.100 113.000 127.200 ;
        RECT 114.200 127.100 114.600 127.200 ;
        RECT 112.200 126.900 114.600 127.100 ;
        RECT 111.000 126.800 111.400 126.900 ;
        RECT 112.600 126.800 114.600 126.900 ;
        RECT 116.600 126.800 117.000 127.200 ;
        RECT 110.200 125.800 110.600 126.600 ;
        RECT 111.100 125.100 111.400 126.800 ;
        RECT 111.800 125.800 112.200 126.600 ;
        RECT 113.400 125.400 113.800 126.200 ;
        RECT 114.200 125.100 114.500 126.800 ;
        RECT 116.700 125.100 117.000 126.800 ;
        RECT 118.200 127.700 118.600 129.900 ;
        RECT 120.300 129.200 120.900 129.900 ;
        RECT 120.300 128.900 121.000 129.200 ;
        RECT 122.600 128.900 123.000 129.900 ;
        RECT 124.800 129.200 125.200 129.900 ;
        RECT 124.800 128.900 125.800 129.200 ;
        RECT 120.600 128.500 121.000 128.900 ;
        RECT 122.700 128.600 123.000 128.900 ;
        RECT 122.700 128.300 124.100 128.600 ;
        RECT 123.700 128.200 124.100 128.300 ;
        RECT 124.600 128.200 125.000 128.600 ;
        RECT 125.400 128.500 125.800 128.900 ;
        RECT 119.700 127.700 120.100 127.800 ;
        RECT 118.200 127.400 120.100 127.700 ;
        RECT 117.400 125.400 117.800 126.200 ;
        RECT 118.200 125.700 118.600 127.400 ;
        RECT 121.700 127.100 122.100 127.200 ;
        RECT 123.800 127.100 124.200 127.200 ;
        RECT 124.600 127.100 124.900 128.200 ;
        RECT 127.000 127.500 127.400 129.900 ;
        RECT 127.800 127.500 128.200 129.900 ;
        RECT 130.000 129.200 130.400 129.900 ;
        RECT 129.400 128.900 130.400 129.200 ;
        RECT 132.200 128.900 132.600 129.900 ;
        RECT 134.300 129.200 134.900 129.900 ;
        RECT 134.200 128.900 134.900 129.200 ;
        RECT 129.400 128.500 129.800 128.900 ;
        RECT 132.200 128.600 132.500 128.900 ;
        RECT 130.200 128.200 130.600 128.600 ;
        RECT 131.100 128.300 132.500 128.600 ;
        RECT 134.200 128.500 134.600 128.900 ;
        RECT 131.100 128.200 131.500 128.300 ;
        RECT 126.200 127.100 127.000 127.200 ;
        RECT 128.200 127.100 129.000 127.200 ;
        RECT 130.300 127.100 130.600 128.200 ;
        RECT 135.100 127.700 135.500 127.800 ;
        RECT 136.600 127.700 137.000 129.900 ;
        RECT 137.400 128.000 137.800 129.900 ;
        RECT 139.000 128.000 139.400 129.900 ;
        RECT 137.400 127.900 139.400 128.000 ;
        RECT 139.800 127.900 140.200 129.900 ;
        RECT 140.900 128.200 141.300 129.900 ;
        RECT 140.900 127.900 141.800 128.200 ;
        RECT 137.500 127.700 139.300 127.900 ;
        RECT 135.100 127.400 137.000 127.700 ;
        RECT 133.100 127.100 133.500 127.200 ;
        RECT 121.500 126.800 133.700 127.100 ;
        RECT 120.600 126.400 121.000 126.500 ;
        RECT 119.100 126.100 121.000 126.400 ;
        RECT 119.100 126.000 119.500 126.100 ;
        RECT 119.900 125.700 120.300 125.800 ;
        RECT 118.200 125.400 120.300 125.700 ;
        RECT 103.000 124.800 103.700 125.100 ;
        RECT 104.000 124.800 104.500 125.100 ;
        RECT 106.200 124.800 106.900 125.100 ;
        RECT 107.200 124.800 107.700 125.100 ;
        RECT 103.400 124.200 103.700 124.800 ;
        RECT 103.400 123.800 103.800 124.200 ;
        RECT 104.100 121.100 104.500 124.800 ;
        RECT 106.600 124.200 106.900 124.800 ;
        RECT 106.600 123.800 107.000 124.200 ;
        RECT 107.300 121.100 107.700 124.800 ;
        RECT 110.700 121.100 111.700 125.100 ;
        RECT 113.700 124.700 114.600 125.100 ;
        RECT 116.600 124.700 117.500 125.100 ;
        RECT 113.700 121.100 114.100 124.700 ;
        RECT 117.100 123.200 117.500 124.700 ;
        RECT 116.600 122.800 117.500 123.200 ;
        RECT 117.100 121.100 117.500 122.800 ;
        RECT 118.200 121.100 118.600 125.400 ;
        RECT 121.500 125.200 121.800 126.800 ;
        RECT 125.100 126.700 125.500 126.800 ;
        RECT 129.700 126.700 130.100 126.800 ;
        RECT 125.900 126.200 126.300 126.300 ;
        RECT 123.800 125.900 126.300 126.200 ;
        RECT 128.900 126.200 129.300 126.300 ;
        RECT 128.900 125.900 131.400 126.200 ;
        RECT 123.800 125.800 124.200 125.900 ;
        RECT 131.000 125.800 131.400 125.900 ;
        RECT 124.600 125.500 127.400 125.600 ;
        RECT 124.500 125.400 127.400 125.500 ;
        RECT 120.600 124.900 121.800 125.200 ;
        RECT 122.500 125.300 127.400 125.400 ;
        RECT 122.500 125.100 124.900 125.300 ;
        RECT 120.600 124.400 120.900 124.900 ;
        RECT 120.200 124.200 120.900 124.400 ;
        RECT 121.700 124.500 122.100 124.600 ;
        RECT 122.500 124.500 122.800 125.100 ;
        RECT 121.700 124.200 122.800 124.500 ;
        RECT 123.100 124.500 125.800 124.800 ;
        RECT 123.100 124.400 123.500 124.500 ;
        RECT 125.400 124.400 125.800 124.500 ;
        RECT 119.800 124.000 120.900 124.200 ;
        RECT 119.800 123.800 120.500 124.000 ;
        RECT 122.300 123.700 122.700 123.800 ;
        RECT 123.700 123.700 124.100 123.800 ;
        RECT 120.600 123.100 121.000 123.500 ;
        RECT 122.300 123.400 124.100 123.700 ;
        RECT 122.700 123.100 123.000 123.400 ;
        RECT 125.400 123.100 125.800 123.500 ;
        RECT 120.300 121.100 120.900 123.100 ;
        RECT 122.600 121.100 123.000 123.100 ;
        RECT 124.800 122.800 125.800 123.100 ;
        RECT 124.800 121.100 125.200 122.800 ;
        RECT 127.000 121.100 127.400 125.300 ;
        RECT 127.800 125.500 130.600 125.600 ;
        RECT 127.800 125.400 130.700 125.500 ;
        RECT 127.800 125.300 132.700 125.400 ;
        RECT 127.800 121.100 128.200 125.300 ;
        RECT 130.300 125.100 132.700 125.300 ;
        RECT 129.400 124.500 132.100 124.800 ;
        RECT 129.400 124.400 129.800 124.500 ;
        RECT 131.700 124.400 132.100 124.500 ;
        RECT 132.400 124.500 132.700 125.100 ;
        RECT 133.400 125.200 133.700 126.800 ;
        RECT 134.200 126.400 134.600 126.500 ;
        RECT 134.200 126.100 136.100 126.400 ;
        RECT 135.700 126.000 136.100 126.100 ;
        RECT 134.900 125.700 135.300 125.800 ;
        RECT 136.600 125.700 137.000 127.400 ;
        RECT 137.800 127.200 138.200 127.400 ;
        RECT 139.800 127.200 140.100 127.900 ;
        RECT 137.400 126.900 138.200 127.200 ;
        RECT 137.400 126.800 137.800 126.900 ;
        RECT 138.900 126.800 140.200 127.200 ;
        RECT 138.200 125.800 138.600 126.600 ;
        RECT 134.900 125.400 137.000 125.700 ;
        RECT 133.400 124.900 134.600 125.200 ;
        RECT 133.100 124.500 133.500 124.600 ;
        RECT 132.400 124.200 133.500 124.500 ;
        RECT 134.300 124.400 134.600 124.900 ;
        RECT 134.300 124.200 135.000 124.400 ;
        RECT 134.300 124.000 135.400 124.200 ;
        RECT 134.700 123.800 135.400 124.000 ;
        RECT 131.100 123.700 131.500 123.800 ;
        RECT 132.500 123.700 132.900 123.800 ;
        RECT 129.400 123.100 129.800 123.500 ;
        RECT 131.100 123.400 132.900 123.700 ;
        RECT 132.200 123.100 132.500 123.400 ;
        RECT 134.200 123.100 134.600 123.500 ;
        RECT 129.400 122.800 130.400 123.100 ;
        RECT 130.000 121.100 130.400 122.800 ;
        RECT 132.200 121.100 132.600 123.100 ;
        RECT 134.300 121.100 134.900 123.100 ;
        RECT 136.600 121.100 137.000 125.400 ;
        RECT 138.900 125.100 139.200 126.800 ;
        RECT 141.400 126.100 141.800 127.900 ;
        RECT 143.000 127.800 143.400 128.600 ;
        RECT 142.200 127.100 142.600 127.600 ;
        RECT 143.000 127.100 143.300 127.800 ;
        RECT 142.200 126.800 143.300 127.100 ;
        RECT 139.800 125.800 141.800 126.100 ;
        RECT 139.800 125.200 140.100 125.800 ;
        RECT 139.800 125.100 140.200 125.200 ;
        RECT 138.700 124.800 139.200 125.100 ;
        RECT 139.500 124.800 140.200 125.100 ;
        RECT 138.700 121.100 139.100 124.800 ;
        RECT 139.500 124.200 139.800 124.800 ;
        RECT 140.600 124.400 141.000 125.200 ;
        RECT 139.400 123.800 139.800 124.200 ;
        RECT 141.400 121.100 141.800 125.800 ;
        RECT 143.800 121.100 144.200 129.900 ;
        RECT 144.600 127.700 145.000 129.900 ;
        RECT 146.700 129.200 147.300 129.900 ;
        RECT 146.700 128.900 147.400 129.200 ;
        RECT 149.000 128.900 149.400 129.900 ;
        RECT 151.200 129.200 151.600 129.900 ;
        RECT 151.200 128.900 152.200 129.200 ;
        RECT 147.000 128.500 147.400 128.900 ;
        RECT 149.100 128.600 149.400 128.900 ;
        RECT 149.100 128.300 150.500 128.600 ;
        RECT 150.100 128.200 150.500 128.300 ;
        RECT 151.000 128.200 151.400 128.600 ;
        RECT 151.800 128.500 152.200 128.900 ;
        RECT 146.100 127.700 146.500 127.800 ;
        RECT 144.600 127.400 146.500 127.700 ;
        RECT 144.600 125.700 145.000 127.400 ;
        RECT 148.100 127.100 148.500 127.200 ;
        RECT 151.000 127.100 151.300 128.200 ;
        RECT 153.400 127.500 153.800 129.900 ;
        RECT 156.600 128.900 157.000 129.900 ;
        RECT 154.200 128.100 154.600 128.200 ;
        RECT 155.800 128.100 156.200 128.600 ;
        RECT 156.700 128.100 157.000 128.900 ;
        RECT 158.300 128.200 158.700 128.600 ;
        RECT 158.200 128.100 158.600 128.200 ;
        RECT 154.200 127.800 156.200 128.100 ;
        RECT 156.600 127.800 158.600 128.100 ;
        RECT 159.000 127.900 159.400 129.900 ;
        RECT 161.500 128.200 161.900 128.600 ;
        RECT 156.700 127.200 157.000 127.800 ;
        RECT 152.600 127.100 153.400 127.200 ;
        RECT 147.900 126.800 153.400 127.100 ;
        RECT 156.600 126.800 157.000 127.200 ;
        RECT 158.200 127.100 158.600 127.200 ;
        RECT 159.100 127.100 159.400 127.900 ;
        RECT 161.400 127.800 161.800 128.200 ;
        RECT 162.200 127.900 162.600 129.900 ;
        RECT 158.200 126.800 159.400 127.100 ;
        RECT 147.000 126.400 147.400 126.500 ;
        RECT 145.500 126.100 147.400 126.400 ;
        RECT 147.900 126.200 148.200 126.800 ;
        RECT 151.500 126.700 151.900 126.800 ;
        RECT 151.000 126.200 151.400 126.300 ;
        RECT 152.300 126.200 152.700 126.300 ;
        RECT 145.500 126.000 145.900 126.100 ;
        RECT 147.800 125.800 148.200 126.200 ;
        RECT 150.200 125.900 152.700 126.200 ;
        RECT 150.200 125.800 150.600 125.900 ;
        RECT 146.300 125.700 146.700 125.800 ;
        RECT 144.600 125.400 146.700 125.700 ;
        RECT 144.600 121.100 145.000 125.400 ;
        RECT 147.900 125.200 148.200 125.800 ;
        RECT 151.000 125.500 153.800 125.600 ;
        RECT 150.900 125.400 153.800 125.500 ;
        RECT 147.000 124.900 148.200 125.200 ;
        RECT 148.900 125.300 153.800 125.400 ;
        RECT 148.900 125.100 151.300 125.300 ;
        RECT 147.000 124.400 147.300 124.900 ;
        RECT 146.600 124.000 147.300 124.400 ;
        RECT 148.100 124.500 148.500 124.600 ;
        RECT 148.900 124.500 149.200 125.100 ;
        RECT 148.100 124.200 149.200 124.500 ;
        RECT 149.500 124.500 152.200 124.800 ;
        RECT 149.500 124.400 149.900 124.500 ;
        RECT 151.800 124.400 152.200 124.500 ;
        RECT 148.700 123.700 149.100 123.800 ;
        RECT 150.100 123.700 150.500 123.800 ;
        RECT 147.000 123.100 147.400 123.500 ;
        RECT 148.700 123.400 150.500 123.700 ;
        RECT 149.100 123.100 149.400 123.400 ;
        RECT 151.800 123.100 152.200 123.500 ;
        RECT 146.700 121.100 147.300 123.100 ;
        RECT 149.000 121.100 149.400 123.100 ;
        RECT 151.200 122.800 152.200 123.100 ;
        RECT 151.200 121.100 151.600 122.800 ;
        RECT 153.400 121.100 153.800 125.300 ;
        RECT 156.700 125.100 157.000 126.800 ;
        RECT 157.400 125.400 157.800 126.200 ;
        RECT 158.200 126.100 158.600 126.200 ;
        RECT 159.100 126.100 159.400 126.800 ;
        RECT 159.800 126.400 160.200 127.200 ;
        RECT 161.400 127.100 161.800 127.200 ;
        RECT 162.300 127.100 162.600 127.900 ;
        RECT 164.600 127.800 165.000 129.900 ;
        RECT 165.400 128.000 165.800 129.900 ;
        RECT 167.000 128.000 167.400 129.900 ;
        RECT 165.400 127.900 167.400 128.000 ;
        RECT 169.400 127.900 169.800 129.900 ;
        RECT 170.100 128.200 170.500 128.600 ;
        RECT 170.200 128.100 170.600 128.200 ;
        RECT 171.000 128.100 171.400 129.900 ;
        RECT 164.700 127.200 165.000 127.800 ;
        RECT 165.500 127.700 167.300 127.900 ;
        RECT 166.600 127.200 167.000 127.400 ;
        RECT 161.400 126.800 162.600 127.100 ;
        RECT 160.600 126.100 161.000 126.200 ;
        RECT 158.200 125.800 159.400 126.100 ;
        RECT 160.200 125.800 161.000 126.100 ;
        RECT 161.400 126.100 161.800 126.200 ;
        RECT 162.300 126.100 162.600 126.800 ;
        RECT 163.000 126.400 163.400 127.200 ;
        RECT 164.600 126.800 165.900 127.200 ;
        RECT 166.600 126.900 167.400 127.200 ;
        RECT 163.800 126.100 164.200 126.200 ;
        RECT 161.400 125.800 162.600 126.100 ;
        RECT 163.400 125.800 164.200 126.100 ;
        RECT 158.300 125.100 158.600 125.800 ;
        RECT 160.200 125.600 160.600 125.800 ;
        RECT 161.500 125.100 161.800 125.800 ;
        RECT 163.400 125.600 163.800 125.800 ;
        RECT 164.600 125.100 165.000 125.200 ;
        RECT 165.600 125.100 165.900 126.800 ;
        RECT 167.000 126.800 167.400 126.900 ;
        RECT 166.200 125.800 166.600 126.600 ;
        RECT 167.000 126.200 167.300 126.800 ;
        RECT 168.600 126.400 169.000 127.200 ;
        RECT 167.000 126.100 167.400 126.200 ;
        RECT 167.800 126.100 168.200 126.200 ;
        RECT 169.400 126.100 169.700 127.900 ;
        RECT 170.200 127.800 171.400 128.100 ;
        RECT 171.800 128.000 172.200 129.900 ;
        RECT 173.400 128.000 173.800 129.900 ;
        RECT 171.800 127.900 173.800 128.000 ;
        RECT 171.100 127.200 171.400 127.800 ;
        RECT 171.900 127.700 173.700 127.900 ;
        RECT 174.200 127.600 174.600 129.900 ;
        RECT 175.800 128.200 176.200 129.900 ;
        RECT 177.700 129.200 178.100 129.900 ;
        RECT 177.400 128.800 178.100 129.200 ;
        RECT 177.700 128.200 178.100 128.800 ;
        RECT 180.100 128.200 180.500 129.900 ;
        RECT 175.800 127.900 176.300 128.200 ;
        RECT 177.700 127.900 178.600 128.200 ;
        RECT 180.100 127.900 181.000 128.200 ;
        RECT 173.000 127.200 173.400 127.400 ;
        RECT 174.200 127.300 175.500 127.600 ;
        RECT 171.000 126.800 172.300 127.200 ;
        RECT 173.000 126.900 173.800 127.200 ;
        RECT 173.400 126.800 173.800 126.900 ;
        RECT 170.200 126.100 170.600 126.200 ;
        RECT 167.000 125.800 168.600 126.100 ;
        RECT 169.400 125.800 170.600 126.100 ;
        RECT 168.200 125.600 168.600 125.800 ;
        RECT 170.200 125.100 170.500 125.800 ;
        RECT 171.000 125.100 171.400 125.200 ;
        RECT 172.000 125.100 172.300 126.800 ;
        RECT 172.600 125.800 173.000 126.600 ;
        RECT 174.300 126.200 174.700 126.600 ;
        RECT 174.200 125.800 174.700 126.200 ;
        RECT 175.200 126.500 175.500 127.300 ;
        RECT 176.000 127.200 176.300 127.900 ;
        RECT 175.800 126.800 176.300 127.200 ;
        RECT 175.200 126.100 175.700 126.500 ;
        RECT 175.200 125.100 175.500 126.100 ;
        RECT 176.000 125.100 176.300 126.800 ;
        RECT 156.600 124.700 157.500 125.100 ;
        RECT 157.100 121.100 157.500 124.700 ;
        RECT 158.200 121.100 158.600 125.100 ;
        RECT 159.000 124.800 161.000 125.100 ;
        RECT 159.000 121.100 159.400 124.800 ;
        RECT 160.600 121.100 161.000 124.800 ;
        RECT 161.400 121.100 161.800 125.100 ;
        RECT 162.200 124.800 164.200 125.100 ;
        RECT 164.600 124.800 165.300 125.100 ;
        RECT 165.600 124.800 166.100 125.100 ;
        RECT 162.200 121.100 162.600 124.800 ;
        RECT 163.800 121.100 164.200 124.800 ;
        RECT 165.000 124.200 165.300 124.800 ;
        RECT 165.000 123.800 165.400 124.200 ;
        RECT 165.700 121.100 166.100 124.800 ;
        RECT 167.800 124.800 169.800 125.100 ;
        RECT 167.800 121.100 168.200 124.800 ;
        RECT 169.400 121.100 169.800 124.800 ;
        RECT 170.200 121.100 170.600 125.100 ;
        RECT 171.000 124.800 171.700 125.100 ;
        RECT 172.000 124.800 172.500 125.100 ;
        RECT 171.400 124.200 171.700 124.800 ;
        RECT 171.400 123.800 171.800 124.200 ;
        RECT 172.100 121.100 172.500 124.800 ;
        RECT 174.200 124.800 175.500 125.100 ;
        RECT 174.200 121.100 174.600 124.800 ;
        RECT 175.800 124.600 176.300 125.100 ;
        RECT 175.800 121.100 176.200 124.600 ;
        RECT 177.400 124.400 177.800 125.200 ;
        RECT 178.200 121.100 178.600 127.900 ;
        RECT 179.800 124.400 180.200 125.200 ;
        RECT 180.600 121.100 181.000 127.900 ;
        RECT 182.200 127.600 182.600 129.900 ;
        RECT 183.800 128.200 184.200 129.900 ;
        RECT 183.800 127.800 184.300 128.200 ;
        RECT 182.200 127.300 183.500 127.600 ;
        RECT 182.300 126.200 182.700 126.600 ;
        RECT 182.200 125.800 182.700 126.200 ;
        RECT 183.200 126.500 183.500 127.300 ;
        RECT 184.000 127.200 184.300 127.800 ;
        RECT 183.800 126.800 184.300 127.200 ;
        RECT 183.200 126.100 183.700 126.500 ;
        RECT 183.200 125.100 183.500 126.100 ;
        RECT 184.000 125.100 184.300 126.800 ;
        RECT 182.200 124.800 183.500 125.100 ;
        RECT 182.200 121.100 182.600 124.800 ;
        RECT 183.800 124.600 184.300 125.100 ;
        RECT 186.200 127.100 186.600 129.900 ;
        RECT 187.000 127.100 187.400 127.200 ;
        RECT 186.200 126.800 187.400 127.100 ;
        RECT 183.800 121.100 184.200 124.600 ;
        RECT 186.200 121.100 186.600 126.800 ;
        RECT 188.600 121.100 189.000 129.900 ;
        RECT 191.000 121.100 191.400 129.900 ;
        RECT 192.600 128.500 193.000 129.500 ;
        RECT 192.600 127.400 192.900 128.500 ;
        RECT 194.700 128.000 195.100 129.500 ;
        RECT 194.700 127.700 195.500 128.000 ;
        RECT 195.100 127.500 195.500 127.700 ;
        RECT 192.600 127.100 194.700 127.400 ;
        RECT 194.200 126.900 194.700 127.100 ;
        RECT 195.200 127.200 195.500 127.500 ;
        RECT 199.000 127.900 199.400 129.900 ;
        RECT 199.700 128.200 200.100 128.600 ;
        RECT 195.200 127.100 196.200 127.200 ;
        RECT 197.400 127.100 197.800 127.200 ;
        RECT 191.800 126.100 192.200 126.200 ;
        RECT 192.600 126.100 193.000 126.600 ;
        RECT 191.800 125.800 193.000 126.100 ;
        RECT 193.400 125.800 193.800 126.600 ;
        RECT 194.200 126.500 194.900 126.900 ;
        RECT 195.200 126.800 197.800 127.100 ;
        RECT 194.200 125.500 194.500 126.500 ;
        RECT 192.600 125.200 194.500 125.500 ;
        RECT 192.600 123.500 192.900 125.200 ;
        RECT 195.200 124.900 195.500 126.800 ;
        RECT 198.200 126.400 198.600 127.200 ;
        RECT 195.800 126.100 196.200 126.200 ;
        RECT 197.400 126.100 197.800 126.200 ;
        RECT 199.000 126.100 199.300 127.900 ;
        RECT 199.800 127.800 200.200 128.200 ;
        RECT 199.800 126.100 200.200 126.200 ;
        RECT 195.800 125.800 198.200 126.100 ;
        RECT 199.000 125.800 200.200 126.100 ;
        RECT 195.800 125.400 196.200 125.800 ;
        RECT 197.800 125.600 198.200 125.800 ;
        RECT 199.800 125.100 200.100 125.800 ;
        RECT 194.700 124.600 195.500 124.900 ;
        RECT 197.400 124.800 199.400 125.100 ;
        RECT 192.600 121.500 193.000 123.500 ;
        RECT 194.700 121.100 195.100 124.600 ;
        RECT 197.400 121.100 197.800 124.800 ;
        RECT 199.000 121.100 199.400 124.800 ;
        RECT 199.800 121.100 200.200 125.100 ;
        RECT 200.600 121.100 201.000 129.900 ;
        RECT 203.000 128.800 203.400 129.900 ;
        RECT 201.400 127.800 201.800 128.600 ;
        RECT 202.200 127.800 202.600 128.600 ;
        RECT 203.100 127.200 203.400 128.800 ;
        RECT 203.000 126.800 203.400 127.200 ;
        RECT 203.100 125.100 203.400 126.800 ;
        RECT 203.800 126.100 204.200 126.200 ;
        RECT 204.600 126.100 205.000 126.200 ;
        RECT 203.800 125.800 205.000 126.100 ;
        RECT 203.800 125.400 204.200 125.800 ;
        RECT 203.000 124.700 203.900 125.100 ;
        RECT 203.500 121.100 203.900 124.700 ;
        RECT 0.600 115.700 1.000 119.900 ;
        RECT 2.800 118.200 3.200 119.900 ;
        RECT 2.200 117.900 3.200 118.200 ;
        RECT 5.000 117.900 5.400 119.900 ;
        RECT 7.100 117.900 7.700 119.900 ;
        RECT 2.200 117.500 2.600 117.900 ;
        RECT 5.000 117.600 5.300 117.900 ;
        RECT 3.900 117.300 5.700 117.600 ;
        RECT 7.000 117.500 7.400 117.900 ;
        RECT 3.900 117.200 4.300 117.300 ;
        RECT 5.300 117.200 5.700 117.300 ;
        RECT 2.200 116.500 2.600 116.600 ;
        RECT 4.500 116.500 4.900 116.600 ;
        RECT 2.200 116.200 4.900 116.500 ;
        RECT 5.200 116.500 6.300 116.800 ;
        RECT 5.200 115.900 5.500 116.500 ;
        RECT 5.900 116.400 6.300 116.500 ;
        RECT 7.100 116.600 7.800 117.000 ;
        RECT 7.100 116.100 7.400 116.600 ;
        RECT 3.100 115.700 5.500 115.900 ;
        RECT 0.600 115.600 5.500 115.700 ;
        RECT 6.200 115.800 7.400 116.100 ;
        RECT 0.600 115.500 3.500 115.600 ;
        RECT 0.600 115.400 3.400 115.500 ;
        RECT 3.800 115.100 4.200 115.200 ;
        RECT 5.400 115.100 5.800 115.200 ;
        RECT 1.700 114.800 5.800 115.100 ;
        RECT 1.700 114.700 2.100 114.800 ;
        RECT 2.500 114.200 2.900 114.300 ;
        RECT 6.200 114.200 6.500 115.800 ;
        RECT 9.400 115.600 9.800 119.900 ;
        RECT 7.700 115.300 9.800 115.600 ;
        RECT 10.200 115.700 10.600 119.900 ;
        RECT 12.400 118.200 12.800 119.900 ;
        RECT 11.800 117.900 12.800 118.200 ;
        RECT 14.600 117.900 15.000 119.900 ;
        RECT 16.700 117.900 17.300 119.900 ;
        RECT 11.800 117.500 12.200 117.900 ;
        RECT 14.600 117.600 14.900 117.900 ;
        RECT 13.500 117.300 15.300 117.600 ;
        RECT 16.600 117.500 17.000 117.900 ;
        RECT 13.500 117.200 13.900 117.300 ;
        RECT 14.900 117.200 15.300 117.300 ;
        RECT 17.100 117.000 17.800 117.200 ;
        RECT 16.700 116.800 17.800 117.000 ;
        RECT 11.800 116.500 12.200 116.600 ;
        RECT 14.100 116.500 14.500 116.600 ;
        RECT 11.800 116.200 14.500 116.500 ;
        RECT 14.800 116.500 15.900 116.800 ;
        RECT 14.800 115.900 15.100 116.500 ;
        RECT 15.500 116.400 15.900 116.500 ;
        RECT 16.700 116.600 17.400 116.800 ;
        RECT 16.700 116.100 17.000 116.600 ;
        RECT 12.700 115.700 15.100 115.900 ;
        RECT 10.200 115.600 15.100 115.700 ;
        RECT 15.800 115.800 17.000 116.100 ;
        RECT 10.200 115.500 13.100 115.600 ;
        RECT 10.200 115.400 13.000 115.500 ;
        RECT 7.700 115.200 8.100 115.300 ;
        RECT 8.500 114.900 8.900 115.000 ;
        RECT 7.000 114.600 8.900 114.900 ;
        RECT 7.000 114.500 7.400 114.600 ;
        RECT 1.000 113.900 6.500 114.200 ;
        RECT 1.000 113.800 1.800 113.900 ;
        RECT 3.000 113.800 3.400 113.900 ;
        RECT 5.900 113.800 6.300 113.900 ;
        RECT 0.600 111.100 1.000 113.500 ;
        RECT 3.100 112.800 3.400 113.800 ;
        RECT 9.400 113.600 9.800 115.300 ;
        RECT 13.400 115.100 13.800 115.200 ;
        RECT 14.200 115.100 14.600 115.200 ;
        RECT 11.300 114.800 14.600 115.100 ;
        RECT 11.300 114.700 11.700 114.800 ;
        RECT 12.100 114.200 12.500 114.300 ;
        RECT 15.800 114.200 16.100 115.800 ;
        RECT 19.000 115.600 19.400 119.900 ;
        RECT 17.300 115.300 19.400 115.600 ;
        RECT 17.300 115.200 17.700 115.300 ;
        RECT 18.100 114.900 18.500 115.000 ;
        RECT 16.600 114.600 18.500 114.900 ;
        RECT 16.600 114.500 17.000 114.600 ;
        RECT 10.600 113.900 16.100 114.200 ;
        RECT 10.600 113.800 11.400 113.900 ;
        RECT 7.900 113.300 9.800 113.600 ;
        RECT 7.900 113.200 8.300 113.300 ;
        RECT 2.200 112.100 2.600 112.500 ;
        RECT 3.000 112.400 3.400 112.800 ;
        RECT 3.900 112.700 4.300 112.800 ;
        RECT 3.900 112.400 5.300 112.700 ;
        RECT 5.000 112.100 5.300 112.400 ;
        RECT 7.000 112.100 7.400 112.500 ;
        RECT 2.200 111.800 3.200 112.100 ;
        RECT 2.800 111.100 3.200 111.800 ;
        RECT 5.000 111.100 5.400 112.100 ;
        RECT 7.000 111.800 7.700 112.100 ;
        RECT 7.100 111.100 7.700 111.800 ;
        RECT 9.400 111.100 9.800 113.300 ;
        RECT 10.200 111.100 10.600 113.500 ;
        RECT 12.700 112.800 13.000 113.900 ;
        RECT 15.500 113.800 15.900 113.900 ;
        RECT 19.000 113.600 19.400 115.300 ;
        RECT 19.800 115.100 20.200 115.200 ;
        RECT 20.600 115.100 21.000 119.900 ;
        RECT 21.400 117.500 21.800 119.500 ;
        RECT 21.400 115.800 21.700 117.500 ;
        RECT 23.500 116.400 23.900 119.900 ;
        RECT 23.500 116.100 24.300 116.400 ;
        RECT 21.400 115.500 23.300 115.800 ;
        RECT 19.800 114.800 21.000 115.100 ;
        RECT 17.500 113.300 19.400 113.600 ;
        RECT 17.500 113.200 17.900 113.300 ;
        RECT 19.000 113.100 19.400 113.300 ;
        RECT 19.800 113.100 20.200 113.200 ;
        RECT 19.000 112.800 20.200 113.100 ;
        RECT 11.800 112.100 12.200 112.500 ;
        RECT 12.600 112.400 13.000 112.800 ;
        RECT 13.500 112.700 13.900 112.800 ;
        RECT 13.500 112.400 14.900 112.700 ;
        RECT 14.600 112.100 14.900 112.400 ;
        RECT 16.600 112.100 17.000 112.500 ;
        RECT 11.800 111.800 12.800 112.100 ;
        RECT 12.400 111.100 12.800 111.800 ;
        RECT 14.600 111.100 15.000 112.100 ;
        RECT 16.600 111.800 17.300 112.100 ;
        RECT 16.700 111.100 17.300 111.800 ;
        RECT 19.000 111.100 19.400 112.800 ;
        RECT 19.800 112.400 20.200 112.800 ;
        RECT 20.600 111.100 21.000 114.800 ;
        RECT 21.400 114.400 21.800 115.200 ;
        RECT 22.200 114.400 22.600 115.200 ;
        RECT 23.000 114.500 23.300 115.500 ;
        RECT 23.000 114.100 23.700 114.500 ;
        RECT 24.000 114.200 24.300 116.100 ;
        RECT 26.200 115.700 26.600 119.900 ;
        RECT 28.400 118.200 28.800 119.900 ;
        RECT 27.800 117.900 28.800 118.200 ;
        RECT 30.600 117.900 31.000 119.900 ;
        RECT 32.700 117.900 33.300 119.900 ;
        RECT 27.800 117.500 28.200 117.900 ;
        RECT 30.600 117.600 30.900 117.900 ;
        RECT 29.500 117.300 31.300 117.600 ;
        RECT 32.600 117.500 33.000 117.900 ;
        RECT 29.500 117.200 29.900 117.300 ;
        RECT 30.900 117.200 31.300 117.300 ;
        RECT 35.000 117.100 35.400 119.900 ;
        RECT 35.800 117.100 36.200 117.200 ;
        RECT 27.800 116.500 28.200 116.600 ;
        RECT 30.100 116.500 30.500 116.600 ;
        RECT 27.800 116.200 30.500 116.500 ;
        RECT 30.800 116.500 31.900 116.800 ;
        RECT 30.800 115.900 31.100 116.500 ;
        RECT 31.500 116.400 31.900 116.500 ;
        RECT 32.700 116.600 33.400 117.000 ;
        RECT 35.000 116.800 36.200 117.100 ;
        RECT 32.700 116.100 33.000 116.600 ;
        RECT 28.700 115.700 31.100 115.900 ;
        RECT 26.200 115.600 31.100 115.700 ;
        RECT 31.800 115.800 33.000 116.100 ;
        RECT 24.600 114.800 25.000 115.600 ;
        RECT 26.200 115.500 29.100 115.600 ;
        RECT 26.200 115.400 29.000 115.500 ;
        RECT 29.400 115.100 29.800 115.200 ;
        RECT 27.300 114.800 29.800 115.100 ;
        RECT 27.300 114.700 27.700 114.800 ;
        RECT 28.100 114.200 28.500 114.300 ;
        RECT 31.800 114.200 32.100 115.800 ;
        RECT 35.000 115.600 35.400 116.800 ;
        RECT 33.300 115.300 35.400 115.600 ;
        RECT 33.300 115.200 33.700 115.300 ;
        RECT 34.100 114.900 34.500 115.000 ;
        RECT 32.600 114.600 34.500 114.900 ;
        RECT 32.600 114.500 33.000 114.600 ;
        RECT 23.000 113.900 23.500 114.100 ;
        RECT 21.400 113.600 23.500 113.900 ;
        RECT 24.000 113.800 25.000 114.200 ;
        RECT 26.600 113.900 32.100 114.200 ;
        RECT 26.600 113.800 27.400 113.900 ;
        RECT 21.400 112.500 21.700 113.600 ;
        RECT 24.000 113.500 24.300 113.800 ;
        RECT 23.900 113.300 24.300 113.500 ;
        RECT 23.500 113.000 24.300 113.300 ;
        RECT 23.500 112.800 24.200 113.000 ;
        RECT 21.400 111.500 21.800 112.500 ;
        RECT 23.500 111.500 23.900 112.800 ;
        RECT 26.200 111.100 26.600 113.500 ;
        RECT 28.700 112.800 29.000 113.900 ;
        RECT 31.500 113.800 31.900 113.900 ;
        RECT 35.000 113.600 35.400 115.300 ;
        RECT 36.600 115.100 37.000 119.900 ;
        RECT 38.600 116.800 39.000 117.200 ;
        RECT 37.400 115.800 37.800 116.600 ;
        RECT 38.600 116.200 38.900 116.800 ;
        RECT 39.300 116.200 39.700 119.900 ;
        RECT 38.200 115.900 38.900 116.200 ;
        RECT 39.200 115.900 39.700 116.200 ;
        RECT 42.700 116.200 43.100 119.900 ;
        RECT 43.400 116.800 43.800 117.200 ;
        RECT 43.500 116.200 43.800 116.800 ;
        RECT 42.700 115.900 43.200 116.200 ;
        RECT 43.500 115.900 44.200 116.200 ;
        RECT 44.600 115.900 45.000 119.900 ;
        RECT 45.400 116.200 45.800 119.900 ;
        RECT 47.000 116.200 47.400 119.900 ;
        RECT 48.600 116.400 49.000 119.900 ;
        RECT 45.400 115.900 47.400 116.200 ;
        RECT 48.500 115.900 49.000 116.400 ;
        RECT 50.200 116.200 50.600 119.900 ;
        RECT 49.300 115.900 50.600 116.200 ;
        RECT 53.900 116.200 54.300 119.900 ;
        RECT 54.600 116.800 55.000 117.200 ;
        RECT 54.700 116.200 55.000 116.800 ;
        RECT 53.900 115.900 54.400 116.200 ;
        RECT 54.700 115.900 55.400 116.200 ;
        RECT 38.200 115.800 38.600 115.900 ;
        RECT 38.200 115.100 38.500 115.800 ;
        RECT 36.600 114.800 38.500 115.100 ;
        RECT 33.500 113.300 35.400 113.600 ;
        RECT 35.800 113.400 36.200 114.200 ;
        RECT 33.500 113.200 33.900 113.300 ;
        RECT 27.800 112.100 28.200 112.500 ;
        RECT 28.600 112.400 29.000 112.800 ;
        RECT 29.500 112.700 29.900 112.800 ;
        RECT 29.500 112.400 30.900 112.700 ;
        RECT 30.600 112.100 30.900 112.400 ;
        RECT 32.600 112.100 33.000 112.500 ;
        RECT 27.800 111.800 28.800 112.100 ;
        RECT 28.400 111.100 28.800 111.800 ;
        RECT 30.600 111.100 31.000 112.100 ;
        RECT 32.600 111.800 33.300 112.100 ;
        RECT 32.700 111.100 33.300 111.800 ;
        RECT 35.000 111.100 35.400 113.300 ;
        RECT 36.600 113.100 37.000 114.800 ;
        RECT 39.200 114.200 39.500 115.900 ;
        RECT 39.800 114.400 40.200 115.200 ;
        RECT 42.200 114.400 42.600 115.200 ;
        RECT 42.900 114.200 43.200 115.900 ;
        RECT 43.800 115.800 44.200 115.900 ;
        RECT 44.700 115.200 45.000 115.900 ;
        RECT 46.600 115.200 47.000 115.400 ;
        RECT 44.600 114.900 45.800 115.200 ;
        RECT 46.600 114.900 47.400 115.200 ;
        RECT 44.600 114.800 45.000 114.900 ;
        RECT 38.200 113.800 39.500 114.200 ;
        RECT 40.600 114.100 41.000 114.200 ;
        RECT 40.200 113.800 41.000 114.100 ;
        RECT 41.400 114.100 41.800 114.200 ;
        RECT 41.400 113.800 42.200 114.100 ;
        RECT 42.900 113.800 44.200 114.200 ;
        RECT 38.300 113.100 38.600 113.800 ;
        RECT 40.200 113.600 40.600 113.800 ;
        RECT 41.800 113.600 42.200 113.800 ;
        RECT 39.100 113.100 40.900 113.300 ;
        RECT 41.500 113.100 43.300 113.300 ;
        RECT 43.800 113.100 44.100 113.800 ;
        RECT 44.600 113.100 45.000 113.200 ;
        RECT 45.500 113.100 45.800 114.900 ;
        RECT 47.000 114.800 47.400 114.900 ;
        RECT 46.200 113.800 46.600 114.600 ;
        RECT 48.500 114.200 48.800 115.900 ;
        RECT 49.300 114.900 49.600 115.900 ;
        RECT 49.100 114.500 49.600 114.900 ;
        RECT 47.800 114.100 48.200 114.200 ;
        RECT 48.500 114.100 49.000 114.200 ;
        RECT 47.800 113.800 49.000 114.100 ;
        RECT 36.600 112.800 37.500 113.100 ;
        RECT 37.100 111.100 37.500 112.800 ;
        RECT 38.200 111.100 38.600 113.100 ;
        RECT 39.000 113.000 41.000 113.100 ;
        RECT 39.000 111.100 39.400 113.000 ;
        RECT 40.600 111.100 41.000 113.000 ;
        RECT 41.400 113.000 43.400 113.100 ;
        RECT 41.400 111.100 41.800 113.000 ;
        RECT 43.000 111.100 43.400 113.000 ;
        RECT 43.800 112.800 45.000 113.100 ;
        RECT 43.800 111.100 44.200 112.800 ;
        RECT 44.700 112.400 45.100 112.800 ;
        RECT 45.400 111.100 45.800 113.100 ;
        RECT 48.500 113.100 48.800 113.800 ;
        RECT 49.300 113.700 49.600 114.500 ;
        RECT 50.100 115.100 50.600 115.200 ;
        RECT 51.000 115.100 51.400 115.200 ;
        RECT 52.600 115.100 53.000 115.200 ;
        RECT 50.100 114.800 53.000 115.100 ;
        RECT 50.100 114.400 50.500 114.800 ;
        RECT 53.400 114.400 53.800 115.200 ;
        RECT 54.100 114.200 54.400 115.900 ;
        RECT 55.000 115.800 55.400 115.900 ;
        RECT 55.800 115.800 56.200 116.600 ;
        RECT 55.000 115.100 55.300 115.800 ;
        RECT 56.600 115.100 57.000 119.900 ;
        RECT 58.200 115.900 58.600 119.900 ;
        RECT 59.000 116.200 59.400 119.900 ;
        RECT 60.600 116.200 61.000 119.900 ;
        RECT 59.000 115.900 61.000 116.200 ;
        RECT 62.700 116.200 63.100 119.900 ;
        RECT 63.400 116.800 63.800 117.200 ;
        RECT 63.500 116.200 63.800 116.800 ;
        RECT 62.700 115.900 63.200 116.200 ;
        RECT 63.500 115.900 64.200 116.200 ;
        RECT 58.300 115.200 58.600 115.900 ;
        RECT 60.200 115.200 60.600 115.400 ;
        RECT 55.000 114.800 57.000 115.100 ;
        RECT 58.200 114.900 59.400 115.200 ;
        RECT 60.200 115.100 61.000 115.200 ;
        RECT 61.400 115.100 61.800 115.200 ;
        RECT 60.200 114.900 61.800 115.100 ;
        RECT 58.200 114.800 58.600 114.900 ;
        RECT 52.600 114.100 53.000 114.200 ;
        RECT 52.600 113.800 53.400 114.100 ;
        RECT 54.100 113.800 55.400 114.200 ;
        RECT 49.300 113.400 50.600 113.700 ;
        RECT 53.000 113.600 53.400 113.800 ;
        RECT 48.500 112.800 49.000 113.100 ;
        RECT 48.600 111.100 49.000 112.800 ;
        RECT 50.200 111.100 50.600 113.400 ;
        RECT 52.700 113.100 54.500 113.300 ;
        RECT 55.000 113.100 55.300 113.800 ;
        RECT 56.600 113.100 57.000 114.800 ;
        RECT 57.400 114.100 57.800 114.200 ;
        RECT 58.200 114.100 58.600 114.200 ;
        RECT 57.400 113.800 58.600 114.100 ;
        RECT 57.400 113.400 57.800 113.800 ;
        RECT 52.600 113.000 54.600 113.100 ;
        RECT 52.600 111.100 53.000 113.000 ;
        RECT 54.200 111.100 54.600 113.000 ;
        RECT 55.000 111.100 55.400 113.100 ;
        RECT 56.100 112.800 57.000 113.100 ;
        RECT 58.200 112.800 58.600 113.200 ;
        RECT 59.100 113.100 59.400 114.900 ;
        RECT 60.600 114.800 61.800 114.900 ;
        RECT 59.800 113.800 60.200 114.600 ;
        RECT 62.200 114.400 62.600 115.200 ;
        RECT 62.900 114.200 63.200 115.900 ;
        RECT 63.800 115.800 64.200 115.900 ;
        RECT 64.600 115.600 65.000 119.900 ;
        RECT 66.700 117.900 67.300 119.900 ;
        RECT 69.000 117.900 69.400 119.900 ;
        RECT 71.200 118.200 71.600 119.900 ;
        RECT 71.200 117.900 72.200 118.200 ;
        RECT 67.000 117.500 67.400 117.900 ;
        RECT 69.100 117.600 69.400 117.900 ;
        RECT 68.700 117.300 70.500 117.600 ;
        RECT 71.800 117.500 72.200 117.900 ;
        RECT 68.700 117.200 69.100 117.300 ;
        RECT 70.100 117.200 70.500 117.300 ;
        RECT 66.600 116.600 67.300 117.000 ;
        RECT 67.000 116.100 67.300 116.600 ;
        RECT 68.100 116.500 69.200 116.800 ;
        RECT 68.100 116.400 68.500 116.500 ;
        RECT 67.000 115.800 68.200 116.100 ;
        RECT 64.600 115.300 66.700 115.600 ;
        RECT 61.400 114.100 61.800 114.200 ;
        RECT 61.400 113.800 62.200 114.100 ;
        RECT 62.900 113.800 64.200 114.200 ;
        RECT 61.800 113.600 62.200 113.800 ;
        RECT 61.500 113.100 63.300 113.300 ;
        RECT 63.800 113.100 64.100 113.800 ;
        RECT 64.600 113.600 65.000 115.300 ;
        RECT 66.300 115.200 66.700 115.300 ;
        RECT 67.900 115.200 68.200 115.800 ;
        RECT 68.900 115.900 69.200 116.500 ;
        RECT 69.500 116.500 69.900 116.600 ;
        RECT 71.800 116.500 72.200 116.600 ;
        RECT 69.500 116.200 72.200 116.500 ;
        RECT 68.900 115.700 71.300 115.900 ;
        RECT 73.400 115.700 73.800 119.900 ;
        RECT 75.000 116.400 75.400 119.900 ;
        RECT 68.900 115.600 73.800 115.700 ;
        RECT 70.900 115.500 73.800 115.600 ;
        RECT 71.000 115.400 73.800 115.500 ;
        RECT 74.900 115.900 75.400 116.400 ;
        RECT 76.600 116.200 77.000 119.900 ;
        RECT 75.700 115.900 77.000 116.200 ;
        RECT 77.400 116.200 77.800 119.900 ;
        RECT 79.000 116.400 79.400 119.900 ;
        RECT 77.400 115.900 78.700 116.200 ;
        RECT 79.000 115.900 79.500 116.400 ;
        RECT 80.600 116.200 81.000 119.900 ;
        RECT 82.200 116.400 82.600 119.900 ;
        RECT 80.600 115.900 81.900 116.200 ;
        RECT 82.200 115.900 82.700 116.400 ;
        RECT 83.800 115.900 84.200 119.900 ;
        RECT 84.600 116.200 85.000 119.900 ;
        RECT 86.200 116.200 86.600 119.900 ;
        RECT 84.600 115.900 86.600 116.200 ;
        RECT 88.300 116.200 88.700 119.900 ;
        RECT 89.000 116.800 89.400 117.200 ;
        RECT 89.100 116.200 89.400 116.800 ;
        RECT 88.300 115.900 88.800 116.200 ;
        RECT 89.100 116.100 89.800 116.200 ;
        RECT 91.000 116.100 91.400 119.900 ;
        RECT 89.100 115.900 91.400 116.100 ;
        RECT 65.500 114.900 65.900 115.000 ;
        RECT 65.500 114.600 67.400 114.900 ;
        RECT 67.800 114.800 68.200 115.200 ;
        RECT 70.200 115.100 70.600 115.200 ;
        RECT 70.200 114.800 72.700 115.100 ;
        RECT 67.000 114.500 67.400 114.600 ;
        RECT 67.900 114.200 68.200 114.800 ;
        RECT 72.300 114.700 72.700 114.800 ;
        RECT 71.500 114.200 71.900 114.300 ;
        RECT 74.900 114.200 75.200 115.900 ;
        RECT 75.700 114.900 76.000 115.900 ;
        RECT 75.500 114.500 76.000 114.900 ;
        RECT 67.900 113.900 73.400 114.200 ;
        RECT 68.100 113.800 68.500 113.900 ;
        RECT 64.600 113.300 66.500 113.600 ;
        RECT 56.100 111.100 56.500 112.800 ;
        RECT 58.300 112.400 58.700 112.800 ;
        RECT 59.000 111.100 59.400 113.100 ;
        RECT 61.400 113.000 63.400 113.100 ;
        RECT 61.400 111.100 61.800 113.000 ;
        RECT 63.000 111.100 63.400 113.000 ;
        RECT 63.800 111.100 64.200 113.100 ;
        RECT 64.600 111.100 65.000 113.300 ;
        RECT 66.100 113.200 66.500 113.300 ;
        RECT 71.000 112.800 71.300 113.900 ;
        RECT 72.600 113.800 73.400 113.900 ;
        RECT 74.200 114.100 74.600 114.200 ;
        RECT 74.900 114.100 75.400 114.200 ;
        RECT 74.200 113.800 75.400 114.100 ;
        RECT 70.100 112.700 70.500 112.800 ;
        RECT 67.000 112.100 67.400 112.500 ;
        RECT 69.100 112.400 70.500 112.700 ;
        RECT 71.000 112.400 71.400 112.800 ;
        RECT 69.100 112.100 69.400 112.400 ;
        RECT 71.800 112.100 72.200 112.500 ;
        RECT 66.700 111.800 67.400 112.100 ;
        RECT 66.700 111.100 67.300 111.800 ;
        RECT 69.000 111.100 69.400 112.100 ;
        RECT 71.200 111.800 72.200 112.100 ;
        RECT 71.200 111.100 71.600 111.800 ;
        RECT 73.400 111.100 73.800 113.500 ;
        RECT 74.900 113.100 75.200 113.800 ;
        RECT 75.700 113.700 76.000 114.500 ;
        RECT 76.500 115.100 77.000 115.200 ;
        RECT 77.400 115.100 77.900 115.200 ;
        RECT 76.500 114.800 77.900 115.100 ;
        RECT 76.500 114.400 76.900 114.800 ;
        RECT 77.500 114.400 77.900 114.800 ;
        RECT 78.400 114.900 78.700 115.900 ;
        RECT 78.400 114.500 78.900 114.900 ;
        RECT 78.400 113.700 78.700 114.500 ;
        RECT 79.200 114.200 79.500 115.900 ;
        RECT 80.600 115.100 81.100 115.200 ;
        RECT 79.000 113.800 79.500 114.200 ;
        RECT 79.800 114.800 81.100 115.100 ;
        RECT 79.800 114.200 80.100 114.800 ;
        RECT 80.700 114.400 81.100 114.800 ;
        RECT 81.600 114.900 81.900 115.900 ;
        RECT 81.600 114.500 82.100 114.900 ;
        RECT 79.800 113.800 80.200 114.200 ;
        RECT 75.700 113.400 77.000 113.700 ;
        RECT 74.900 112.800 75.400 113.100 ;
        RECT 75.000 111.100 75.400 112.800 ;
        RECT 76.600 111.100 77.000 113.400 ;
        RECT 77.400 113.400 78.700 113.700 ;
        RECT 77.400 111.100 77.800 113.400 ;
        RECT 79.200 113.100 79.500 113.800 ;
        RECT 81.600 113.700 81.900 114.500 ;
        RECT 82.400 114.200 82.700 115.900 ;
        RECT 83.900 115.200 84.200 115.900 ;
        RECT 85.800 115.200 86.200 115.400 ;
        RECT 83.800 114.900 85.000 115.200 ;
        RECT 85.800 115.100 86.600 115.200 ;
        RECT 87.000 115.100 87.400 115.200 ;
        RECT 85.800 114.900 87.400 115.100 ;
        RECT 83.800 114.800 84.200 114.900 ;
        RECT 82.200 113.800 82.700 114.200 ;
        RECT 83.000 114.100 83.400 114.200 ;
        RECT 84.700 114.100 85.000 114.900 ;
        RECT 86.200 114.800 87.400 114.900 ;
        RECT 83.000 113.800 85.000 114.100 ;
        RECT 85.400 113.800 85.800 114.600 ;
        RECT 87.800 114.400 88.200 115.200 ;
        RECT 88.500 114.200 88.800 115.900 ;
        RECT 89.400 115.800 91.400 115.900 ;
        RECT 91.800 115.800 92.200 116.600 ;
        RECT 86.200 114.100 86.600 114.200 ;
        RECT 87.000 114.100 87.400 114.200 ;
        RECT 86.200 113.800 87.800 114.100 ;
        RECT 88.500 113.800 89.800 114.200 ;
        RECT 79.000 112.800 79.500 113.100 ;
        RECT 80.600 113.400 81.900 113.700 ;
        RECT 79.000 111.100 79.400 112.800 ;
        RECT 80.600 111.100 81.000 113.400 ;
        RECT 82.400 113.100 82.700 113.800 ;
        RECT 82.200 112.800 82.700 113.100 ;
        RECT 83.800 112.800 84.200 113.200 ;
        RECT 84.700 113.100 85.000 113.800 ;
        RECT 87.400 113.600 87.800 113.800 ;
        RECT 87.100 113.100 88.900 113.300 ;
        RECT 89.400 113.100 89.700 113.800 ;
        RECT 90.200 113.400 90.600 114.200 ;
        RECT 91.000 113.100 91.400 115.800 ;
        RECT 92.600 115.700 93.000 119.900 ;
        RECT 94.800 118.200 95.200 119.900 ;
        RECT 94.200 117.900 95.200 118.200 ;
        RECT 97.000 117.900 97.400 119.900 ;
        RECT 99.100 117.900 99.700 119.900 ;
        RECT 94.200 117.500 94.600 117.900 ;
        RECT 97.000 117.600 97.300 117.900 ;
        RECT 95.900 117.300 97.700 117.600 ;
        RECT 99.000 117.500 99.400 117.900 ;
        RECT 95.900 117.200 96.300 117.300 ;
        RECT 97.300 117.200 97.700 117.300 ;
        RECT 94.200 116.500 94.600 116.600 ;
        RECT 96.500 116.500 96.900 116.600 ;
        RECT 94.200 116.200 96.900 116.500 ;
        RECT 97.200 116.500 98.300 116.800 ;
        RECT 97.200 115.900 97.500 116.500 ;
        RECT 97.900 116.400 98.300 116.500 ;
        RECT 99.100 116.600 99.800 117.000 ;
        RECT 99.100 116.100 99.400 116.600 ;
        RECT 95.100 115.700 97.500 115.900 ;
        RECT 92.600 115.600 97.500 115.700 ;
        RECT 98.200 115.800 99.400 116.100 ;
        RECT 92.600 115.500 95.500 115.600 ;
        RECT 92.600 115.400 95.400 115.500 ;
        RECT 95.800 115.100 96.200 115.200 ;
        RECT 96.600 115.100 97.000 115.200 ;
        RECT 93.700 114.800 97.000 115.100 ;
        RECT 93.700 114.700 94.100 114.800 ;
        RECT 94.500 114.200 94.900 114.300 ;
        RECT 98.200 114.200 98.500 115.800 ;
        RECT 101.400 115.600 101.800 119.900 ;
        RECT 99.700 115.300 101.800 115.600 ;
        RECT 99.700 115.200 100.100 115.300 ;
        RECT 100.500 114.900 100.900 115.000 ;
        RECT 99.000 114.600 100.900 114.900 ;
        RECT 99.000 114.500 99.400 114.600 ;
        RECT 93.000 113.900 98.500 114.200 ;
        RECT 93.000 113.800 93.800 113.900 ;
        RECT 82.200 111.100 82.600 112.800 ;
        RECT 83.900 112.400 84.300 112.800 ;
        RECT 84.600 111.100 85.000 113.100 ;
        RECT 87.000 113.000 89.000 113.100 ;
        RECT 87.000 111.100 87.400 113.000 ;
        RECT 88.600 111.100 89.000 113.000 ;
        RECT 89.400 111.100 89.800 113.100 ;
        RECT 91.000 112.800 91.900 113.100 ;
        RECT 91.500 111.100 91.900 112.800 ;
        RECT 92.600 111.100 93.000 113.500 ;
        RECT 95.100 112.800 95.400 113.900 ;
        RECT 97.900 113.800 98.300 113.900 ;
        RECT 101.400 113.600 101.800 115.300 ;
        RECT 104.600 115.100 105.000 119.900 ;
        RECT 106.600 116.800 107.000 117.200 ;
        RECT 105.400 115.800 105.800 116.600 ;
        RECT 106.600 116.200 106.900 116.800 ;
        RECT 107.300 116.200 107.700 119.900 ;
        RECT 106.200 115.900 106.900 116.200 ;
        RECT 107.200 115.900 107.700 116.200 ;
        RECT 109.400 116.200 109.800 119.900 ;
        RECT 111.000 116.400 111.400 119.900 ;
        RECT 109.400 115.900 110.700 116.200 ;
        RECT 111.000 115.900 111.500 116.400 ;
        RECT 112.600 116.200 113.000 119.900 ;
        RECT 114.800 119.200 115.600 119.900 ;
        RECT 114.200 118.800 115.600 119.200 ;
        RECT 113.400 116.200 113.800 116.300 ;
        RECT 114.800 116.200 115.600 118.800 ;
        RECT 112.600 115.900 113.800 116.200 ;
        RECT 114.600 115.900 115.600 116.200 ;
        RECT 116.700 116.200 117.100 116.300 ;
        RECT 117.400 116.200 117.800 119.900 ;
        RECT 119.000 116.400 119.400 119.900 ;
        RECT 116.700 115.900 117.800 116.200 ;
        RECT 106.200 115.800 106.600 115.900 ;
        RECT 106.200 115.100 106.500 115.800 ;
        RECT 104.600 114.800 106.500 115.100 ;
        RECT 102.200 114.100 102.600 114.200 ;
        RECT 103.800 114.100 104.200 114.200 ;
        RECT 102.200 113.800 104.200 114.100 ;
        RECT 99.900 113.300 101.800 113.600 ;
        RECT 103.800 113.400 104.200 113.800 ;
        RECT 99.900 113.200 100.300 113.300 ;
        RECT 94.200 112.100 94.600 112.500 ;
        RECT 95.000 112.400 95.400 112.800 ;
        RECT 95.900 112.700 96.300 112.800 ;
        RECT 95.900 112.400 97.300 112.700 ;
        RECT 97.000 112.100 97.300 112.400 ;
        RECT 99.000 112.100 99.400 112.500 ;
        RECT 101.400 112.100 101.800 113.300 ;
        RECT 104.600 113.100 105.000 114.800 ;
        RECT 107.200 114.200 107.500 115.900 ;
        RECT 107.800 114.400 108.200 115.200 ;
        RECT 109.400 114.800 109.900 115.200 ;
        RECT 109.500 114.400 109.900 114.800 ;
        RECT 110.400 114.900 110.700 115.900 ;
        RECT 110.400 114.500 110.900 114.900 ;
        RECT 106.200 113.800 107.500 114.200 ;
        RECT 108.600 114.100 109.000 114.200 ;
        RECT 108.200 113.800 109.000 114.100 ;
        RECT 106.300 113.100 106.600 113.800 ;
        RECT 108.200 113.600 108.600 113.800 ;
        RECT 110.400 113.700 110.700 114.500 ;
        RECT 111.200 114.200 111.500 115.900 ;
        RECT 114.600 115.200 114.900 115.900 ;
        RECT 116.700 115.600 117.000 115.900 ;
        RECT 115.300 115.300 117.000 115.600 ;
        RECT 118.900 115.800 119.400 116.400 ;
        RECT 120.600 116.200 121.000 119.900 ;
        RECT 122.500 119.200 122.900 119.900 ;
        RECT 122.500 118.800 123.400 119.200 ;
        RECT 121.800 116.800 122.200 117.200 ;
        RECT 121.800 116.200 122.100 116.800 ;
        RECT 122.500 116.200 122.900 118.800 ;
        RECT 119.700 115.900 121.000 116.200 ;
        RECT 121.400 115.900 122.100 116.200 ;
        RECT 122.400 115.900 122.900 116.200 ;
        RECT 124.600 116.200 125.000 119.900 ;
        RECT 126.200 116.200 126.600 119.900 ;
        RECT 124.600 115.900 126.600 116.200 ;
        RECT 127.000 116.100 127.400 119.900 ;
        RECT 128.900 118.200 129.300 119.900 ;
        RECT 128.900 117.800 129.800 118.200 ;
        RECT 128.200 116.800 128.600 117.200 ;
        RECT 128.200 116.200 128.500 116.800 ;
        RECT 128.900 116.200 129.300 117.800 ;
        RECT 127.800 116.100 128.500 116.200 ;
        RECT 127.000 115.900 128.500 116.100 ;
        RECT 128.800 115.900 129.300 116.200 ;
        RECT 115.300 115.200 115.700 115.300 ;
        RECT 114.200 114.900 114.900 115.200 ;
        RECT 116.400 114.900 116.800 115.000 ;
        RECT 114.200 114.800 115.100 114.900 ;
        RECT 114.600 114.600 115.100 114.800 ;
        RECT 111.000 114.100 111.500 114.200 ;
        RECT 111.800 114.100 112.200 114.200 ;
        RECT 111.000 113.800 112.200 114.100 ;
        RECT 112.600 113.800 113.400 114.200 ;
        RECT 114.000 113.800 114.400 114.200 ;
        RECT 109.400 113.400 110.700 113.700 ;
        RECT 107.100 113.100 108.900 113.300 ;
        RECT 104.600 112.800 105.500 113.100 ;
        RECT 102.200 112.100 102.600 112.200 ;
        RECT 94.200 111.800 95.200 112.100 ;
        RECT 94.800 111.100 95.200 111.800 ;
        RECT 97.000 111.100 97.400 112.100 ;
        RECT 99.000 111.800 99.700 112.100 ;
        RECT 99.100 111.100 99.700 111.800 ;
        RECT 101.400 111.800 102.600 112.100 ;
        RECT 101.400 111.100 101.800 111.800 ;
        RECT 105.100 111.100 105.500 112.800 ;
        RECT 106.200 111.100 106.600 113.100 ;
        RECT 107.000 113.000 109.000 113.100 ;
        RECT 107.000 111.100 107.400 113.000 ;
        RECT 108.600 111.100 109.000 113.000 ;
        RECT 109.400 111.100 109.800 113.400 ;
        RECT 111.200 113.100 111.500 113.800 ;
        RECT 114.100 113.600 114.400 113.800 ;
        RECT 113.400 113.400 113.800 113.500 ;
        RECT 111.000 112.800 111.500 113.100 ;
        RECT 112.600 113.100 113.800 113.400 ;
        RECT 114.100 113.200 114.500 113.600 ;
        RECT 111.000 111.100 111.400 112.800 ;
        RECT 112.600 111.100 113.000 113.100 ;
        RECT 114.800 112.900 115.100 114.600 ;
        RECT 115.500 114.600 116.800 114.900 ;
        RECT 115.500 114.300 115.800 114.600 ;
        RECT 115.400 113.900 115.800 114.300 ;
        RECT 118.900 114.200 119.200 115.800 ;
        RECT 119.700 114.900 120.000 115.900 ;
        RECT 121.400 115.800 121.800 115.900 ;
        RECT 119.500 114.500 120.000 114.900 ;
        RECT 117.000 114.100 117.800 114.200 ;
        RECT 116.100 113.800 117.800 114.100 ;
        RECT 118.900 113.800 119.400 114.200 ;
        RECT 116.100 113.600 116.400 113.800 ;
        RECT 115.400 113.300 116.400 113.600 ;
        RECT 116.700 113.400 117.100 113.500 ;
        RECT 115.400 113.200 116.200 113.300 ;
        RECT 116.700 113.100 117.800 113.400 ;
        RECT 114.800 111.100 115.600 112.900 ;
        RECT 117.400 111.100 117.800 113.100 ;
        RECT 118.900 113.100 119.200 113.800 ;
        RECT 119.700 113.700 120.000 114.500 ;
        RECT 120.500 114.800 121.000 115.200 ;
        RECT 120.500 114.400 120.900 114.800 ;
        RECT 122.400 114.200 122.700 115.900 ;
        RECT 127.000 115.800 128.200 115.900 ;
        RECT 125.000 115.200 125.400 115.400 ;
        RECT 127.000 115.200 127.300 115.800 ;
        RECT 123.000 115.100 123.400 115.200 ;
        RECT 123.800 115.100 124.200 115.200 ;
        RECT 123.000 114.800 124.200 115.100 ;
        RECT 124.600 114.900 125.400 115.200 ;
        RECT 126.200 114.900 127.400 115.200 ;
        RECT 124.600 114.800 125.000 114.900 ;
        RECT 123.000 114.400 123.400 114.800 ;
        RECT 121.400 113.800 122.700 114.200 ;
        RECT 123.800 114.100 124.200 114.200 ;
        RECT 123.400 113.800 124.200 114.100 ;
        RECT 125.400 113.800 125.800 114.600 ;
        RECT 119.700 113.400 121.000 113.700 ;
        RECT 118.900 112.800 119.400 113.100 ;
        RECT 119.000 111.100 119.400 112.800 ;
        RECT 120.600 111.100 121.000 113.400 ;
        RECT 121.500 113.100 121.800 113.800 ;
        RECT 123.400 113.600 123.800 113.800 ;
        RECT 122.300 113.100 124.100 113.300 ;
        RECT 126.200 113.100 126.500 114.900 ;
        RECT 127.000 114.800 127.400 114.900 ;
        RECT 128.800 114.200 129.100 115.900 ;
        RECT 129.400 114.400 129.800 115.200 ;
        RECT 127.800 113.800 129.100 114.200 ;
        RECT 130.200 114.100 130.600 114.200 ;
        RECT 129.800 113.800 130.600 114.100 ;
        RECT 121.400 111.100 121.800 113.100 ;
        RECT 122.200 113.000 124.200 113.100 ;
        RECT 122.200 111.100 122.600 113.000 ;
        RECT 123.800 111.100 124.200 113.000 ;
        RECT 126.200 111.100 126.600 113.100 ;
        RECT 127.000 112.800 127.400 113.200 ;
        RECT 127.900 113.100 128.200 113.800 ;
        RECT 129.800 113.600 130.200 113.800 ;
        RECT 131.000 113.400 131.400 114.200 ;
        RECT 131.800 114.100 132.200 119.900 ;
        RECT 132.600 115.800 133.000 116.600 ;
        RECT 134.200 116.000 134.600 119.900 ;
        RECT 135.800 117.600 136.200 119.900 ;
        RECT 134.100 115.600 134.600 116.000 ;
        RECT 134.900 117.300 136.200 117.600 ;
        RECT 134.900 116.500 135.200 117.300 ;
        RECT 137.400 117.200 137.800 119.900 ;
        RECT 139.000 118.500 139.400 119.900 ;
        RECT 139.800 118.500 140.200 119.900 ;
        RECT 140.600 118.500 141.000 119.900 ;
        RECT 138.100 117.200 140.200 117.600 ;
        RECT 136.500 116.800 137.800 117.200 ;
        RECT 141.400 116.800 141.800 119.900 ;
        RECT 143.000 117.500 143.400 119.900 ;
        RECT 144.600 117.500 145.000 119.900 ;
        RECT 145.400 118.500 145.800 119.900 ;
        RECT 146.200 118.500 146.600 119.900 ;
        RECT 147.800 117.600 148.200 119.900 ;
        RECT 149.400 118.200 149.800 119.900 ;
        RECT 149.400 117.900 149.900 118.200 ;
        RECT 149.600 117.600 149.900 117.900 ;
        RECT 147.200 117.200 149.300 117.600 ;
        RECT 149.600 117.300 150.600 117.600 ;
        RECT 143.000 116.800 144.300 117.200 ;
        RECT 144.600 116.900 147.500 117.200 ;
        RECT 149.000 117.000 149.300 117.200 ;
        RECT 139.000 116.500 139.400 116.600 ;
        RECT 134.900 116.200 139.400 116.500 ;
        RECT 140.600 116.500 141.000 116.600 ;
        RECT 144.600 116.500 144.900 116.900 ;
        RECT 147.800 116.600 148.500 116.900 ;
        RECT 149.000 116.600 149.800 117.000 ;
        RECT 140.600 116.200 144.900 116.500 ;
        RECT 145.400 116.500 148.500 116.600 ;
        RECT 145.400 116.300 148.100 116.500 ;
        RECT 145.400 116.200 145.800 116.300 ;
        RECT 132.600 114.100 133.000 114.200 ;
        RECT 131.800 113.800 133.000 114.100 ;
        RECT 128.700 113.100 130.500 113.300 ;
        RECT 131.800 113.100 132.200 113.800 ;
        RECT 134.100 113.400 134.500 115.600 ;
        RECT 134.900 115.300 135.200 116.200 ;
        RECT 134.800 115.000 135.200 115.300 ;
        RECT 138.200 115.000 149.900 115.300 ;
        RECT 134.800 114.000 135.100 115.000 ;
        RECT 138.200 114.700 138.600 115.000 ;
        RECT 147.000 114.800 147.400 115.000 ;
        RECT 149.400 114.900 149.900 115.000 ;
        RECT 149.400 114.800 149.800 114.900 ;
        RECT 135.400 114.300 137.300 114.700 ;
        RECT 134.800 113.700 135.400 114.000 ;
        RECT 126.900 112.400 127.300 112.800 ;
        RECT 127.800 111.100 128.200 113.100 ;
        RECT 128.600 113.000 130.600 113.100 ;
        RECT 128.600 111.100 129.000 113.000 ;
        RECT 130.200 111.100 130.600 113.000 ;
        RECT 131.800 112.800 132.700 113.100 ;
        RECT 134.100 113.000 134.600 113.400 ;
        RECT 132.300 111.100 132.700 112.800 ;
        RECT 134.200 111.100 134.600 113.000 ;
        RECT 135.000 111.100 135.400 113.700 ;
        RECT 136.900 113.700 137.300 114.300 ;
        RECT 136.900 113.400 137.800 113.700 ;
        RECT 137.400 113.100 137.800 113.400 ;
        RECT 139.800 113.200 140.200 114.600 ;
        RECT 141.400 114.300 143.000 114.700 ;
        RECT 144.900 114.300 145.900 114.700 ;
        RECT 150.200 114.500 150.600 117.300 ;
        RECT 151.300 116.300 151.700 119.900 ;
        RECT 151.300 115.900 152.200 116.300 ;
        RECT 155.000 115.900 155.400 119.900 ;
        RECT 155.800 116.200 156.200 119.900 ;
        RECT 157.400 116.200 157.800 119.900 ;
        RECT 155.800 115.900 157.800 116.200 ;
        RECT 158.200 115.900 158.600 119.900 ;
        RECT 159.000 116.200 159.400 119.900 ;
        RECT 160.600 116.200 161.000 119.900 ;
        RECT 161.400 117.900 161.800 119.900 ;
        RECT 161.500 117.800 161.800 117.900 ;
        RECT 163.000 117.900 163.400 119.900 ;
        RECT 165.900 119.200 166.300 119.900 ;
        RECT 165.400 118.800 166.300 119.200 ;
        RECT 163.000 117.800 163.300 117.900 ;
        RECT 161.500 117.500 163.300 117.800 ;
        RECT 161.500 116.200 161.800 117.500 ;
        RECT 162.200 116.400 162.600 117.200 ;
        RECT 165.900 116.200 166.300 118.800 ;
        RECT 168.600 118.200 169.000 119.900 ;
        RECT 168.500 117.900 169.000 118.200 ;
        RECT 168.500 117.600 168.800 117.900 ;
        RECT 170.200 117.600 170.600 119.900 ;
        RECT 171.800 118.500 172.200 119.900 ;
        RECT 172.600 118.500 173.000 119.900 ;
        RECT 167.800 117.300 168.800 117.600 ;
        RECT 166.600 116.800 167.000 117.200 ;
        RECT 166.700 116.200 167.000 116.800 ;
        RECT 159.000 115.900 161.000 116.200 ;
        RECT 151.800 115.800 152.200 115.900 ;
        RECT 151.000 114.800 151.400 115.600 ;
        RECT 141.200 113.900 141.600 114.000 ;
        RECT 141.200 113.600 143.400 113.900 ;
        RECT 143.000 113.500 143.400 113.600 ;
        RECT 143.800 113.400 144.200 114.200 ;
        RECT 137.400 112.700 138.600 113.100 ;
        RECT 139.800 112.800 140.300 113.200 ;
        RECT 141.800 112.800 142.600 113.200 ;
        RECT 143.000 113.100 143.400 113.200 ;
        RECT 144.900 113.100 145.300 114.300 ;
        RECT 146.200 114.100 150.600 114.500 ;
        RECT 147.900 113.400 149.400 113.800 ;
        RECT 147.900 113.100 148.300 113.400 ;
        RECT 143.000 112.800 145.300 113.100 ;
        RECT 138.200 111.100 138.600 112.700 ;
        RECT 147.000 112.700 148.300 113.100 ;
        RECT 139.000 111.100 139.400 112.500 ;
        RECT 139.800 111.100 140.200 112.500 ;
        RECT 140.600 111.100 141.000 112.500 ;
        RECT 141.400 111.100 141.800 112.500 ;
        RECT 143.000 111.100 143.400 112.500 ;
        RECT 144.600 111.100 145.000 112.500 ;
        RECT 145.400 111.100 145.800 112.500 ;
        RECT 146.200 111.100 146.600 112.500 ;
        RECT 147.000 111.100 147.400 112.700 ;
        RECT 150.200 111.100 150.600 114.100 ;
        RECT 151.800 114.200 152.100 115.800 ;
        RECT 155.100 115.200 155.400 115.900 ;
        RECT 157.000 115.200 157.400 115.400 ;
        RECT 158.300 115.200 158.600 115.900 ;
        RECT 161.400 115.800 161.800 116.200 ;
        RECT 160.200 115.200 160.600 115.400 ;
        RECT 155.000 114.900 156.200 115.200 ;
        RECT 157.000 114.900 157.800 115.200 ;
        RECT 155.000 114.800 155.400 114.900 ;
        RECT 151.800 113.800 152.200 114.200 ;
        RECT 151.800 112.100 152.100 113.800 ;
        RECT 152.600 112.400 153.000 113.200 ;
        RECT 154.200 113.100 154.600 113.200 ;
        RECT 155.000 113.100 155.400 113.200 ;
        RECT 155.900 113.100 156.200 114.900 ;
        RECT 157.400 114.800 157.800 114.900 ;
        RECT 158.200 114.900 159.400 115.200 ;
        RECT 160.200 114.900 161.000 115.200 ;
        RECT 158.200 114.800 158.600 114.900 ;
        RECT 156.600 113.800 157.000 114.600 ;
        RECT 159.100 113.200 159.400 114.900 ;
        RECT 160.600 114.800 161.000 114.900 ;
        RECT 159.800 113.800 160.200 114.600 ;
        RECT 161.500 114.200 161.800 115.800 ;
        RECT 163.800 115.400 164.200 116.200 ;
        RECT 165.900 115.900 166.400 116.200 ;
        RECT 166.700 115.900 167.400 116.200 ;
        RECT 162.600 114.800 163.400 115.200 ;
        RECT 165.400 114.400 165.800 115.200 ;
        RECT 166.100 114.200 166.400 115.900 ;
        RECT 167.000 115.800 167.400 115.900 ;
        RECT 167.800 114.500 168.200 117.300 ;
        RECT 169.100 117.200 171.200 117.600 ;
        RECT 173.400 117.500 173.800 119.900 ;
        RECT 175.000 117.500 175.400 119.900 ;
        RECT 169.100 117.000 169.400 117.200 ;
        RECT 168.600 116.600 169.400 117.000 ;
        RECT 170.900 116.900 173.800 117.200 ;
        RECT 169.900 116.600 170.600 116.900 ;
        RECT 169.900 116.500 173.000 116.600 ;
        RECT 170.300 116.300 173.000 116.500 ;
        RECT 172.600 116.200 173.000 116.300 ;
        RECT 173.500 116.500 173.800 116.900 ;
        RECT 174.100 116.800 175.400 117.200 ;
        RECT 176.600 116.800 177.000 119.900 ;
        RECT 177.400 118.500 177.800 119.900 ;
        RECT 178.200 118.500 178.600 119.900 ;
        RECT 179.000 118.500 179.400 119.900 ;
        RECT 178.200 117.200 180.300 117.600 ;
        RECT 180.600 117.200 181.000 119.900 ;
        RECT 182.200 117.600 182.600 119.900 ;
        RECT 182.200 117.300 183.500 117.600 ;
        RECT 180.600 116.800 181.900 117.200 ;
        RECT 177.400 116.500 177.800 116.600 ;
        RECT 173.500 116.200 177.800 116.500 ;
        RECT 179.000 116.500 179.400 116.600 ;
        RECT 183.200 116.500 183.500 117.300 ;
        RECT 179.000 116.200 183.500 116.500 ;
        RECT 183.200 115.300 183.500 116.200 ;
        RECT 183.800 116.000 184.200 119.900 ;
        RECT 183.800 115.600 184.300 116.000 ;
        RECT 168.500 115.000 180.200 115.300 ;
        RECT 183.200 115.000 183.600 115.300 ;
        RECT 168.500 114.900 168.900 115.000 ;
        RECT 169.400 114.800 169.800 115.000 ;
        RECT 171.000 114.800 171.400 115.000 ;
        RECT 179.800 114.700 180.200 115.000 ;
        RECT 161.500 114.100 162.300 114.200 ;
        RECT 164.600 114.100 165.000 114.200 ;
        RECT 161.500 113.900 162.400 114.100 ;
        RECT 154.200 112.800 155.400 113.100 ;
        RECT 155.100 112.400 155.500 112.800 ;
        RECT 151.800 111.100 152.200 112.100 ;
        RECT 155.800 111.100 156.200 113.100 ;
        RECT 158.200 112.800 158.600 113.200 ;
        RECT 158.300 112.400 158.700 112.800 ;
        RECT 159.000 111.100 159.400 113.200 ;
        RECT 162.000 111.100 162.400 113.900 ;
        RECT 164.600 113.800 165.400 114.100 ;
        RECT 166.100 113.800 167.400 114.200 ;
        RECT 167.800 114.100 172.200 114.500 ;
        RECT 172.500 114.300 173.500 114.700 ;
        RECT 175.400 114.300 177.000 114.700 ;
        RECT 165.000 113.600 165.400 113.800 ;
        RECT 164.700 113.100 166.500 113.300 ;
        RECT 167.000 113.100 167.300 113.800 ;
        RECT 164.600 113.000 166.600 113.100 ;
        RECT 164.600 111.100 165.000 113.000 ;
        RECT 166.200 111.100 166.600 113.000 ;
        RECT 167.000 111.100 167.400 113.100 ;
        RECT 167.800 111.100 168.200 114.100 ;
        RECT 169.000 113.400 170.500 113.800 ;
        RECT 170.100 113.100 170.500 113.400 ;
        RECT 173.100 113.100 173.500 114.300 ;
        RECT 174.200 113.400 174.600 114.200 ;
        RECT 176.800 113.900 177.200 114.000 ;
        RECT 175.000 113.600 177.200 113.900 ;
        RECT 175.000 113.500 175.400 113.600 ;
        RECT 178.200 113.200 178.600 114.600 ;
        RECT 181.100 114.300 183.000 114.700 ;
        RECT 181.100 113.700 181.500 114.300 ;
        RECT 183.300 114.000 183.600 115.000 ;
        RECT 175.000 113.100 175.400 113.200 ;
        RECT 170.100 112.700 171.400 113.100 ;
        RECT 173.100 112.800 175.400 113.100 ;
        RECT 175.800 112.800 176.600 113.200 ;
        RECT 178.100 112.800 178.600 113.200 ;
        RECT 180.600 113.400 181.500 113.700 ;
        RECT 183.000 113.700 183.600 114.000 ;
        RECT 180.600 113.100 181.000 113.400 ;
        RECT 171.000 111.100 171.400 112.700 ;
        RECT 179.800 112.700 181.000 113.100 ;
        RECT 171.800 111.100 172.200 112.500 ;
        RECT 172.600 111.100 173.000 112.500 ;
        RECT 173.400 111.100 173.800 112.500 ;
        RECT 175.000 111.100 175.400 112.500 ;
        RECT 176.600 111.100 177.000 112.500 ;
        RECT 177.400 111.100 177.800 112.500 ;
        RECT 178.200 111.100 178.600 112.500 ;
        RECT 179.000 111.100 179.400 112.500 ;
        RECT 179.800 111.100 180.200 112.700 ;
        RECT 183.000 111.100 183.400 113.700 ;
        RECT 183.900 113.400 184.300 115.600 ;
        RECT 183.800 113.000 184.300 113.400 ;
        RECT 185.400 115.600 185.800 119.900 ;
        RECT 187.500 117.900 188.100 119.900 ;
        RECT 189.800 117.900 190.200 119.900 ;
        RECT 192.000 118.200 192.400 119.900 ;
        RECT 192.000 117.900 193.000 118.200 ;
        RECT 187.800 117.500 188.200 117.900 ;
        RECT 189.900 117.600 190.200 117.900 ;
        RECT 189.500 117.300 191.300 117.600 ;
        RECT 192.600 117.500 193.000 117.900 ;
        RECT 189.500 117.200 189.900 117.300 ;
        RECT 190.900 117.200 191.300 117.300 ;
        RECT 187.400 116.600 188.100 117.000 ;
        RECT 187.800 116.100 188.100 116.600 ;
        RECT 188.900 116.500 190.000 116.800 ;
        RECT 188.900 116.400 189.300 116.500 ;
        RECT 187.800 115.800 189.000 116.100 ;
        RECT 185.400 115.300 187.500 115.600 ;
        RECT 185.400 113.600 185.800 115.300 ;
        RECT 187.100 115.200 187.500 115.300 ;
        RECT 188.700 115.200 189.000 115.800 ;
        RECT 189.700 115.900 190.000 116.500 ;
        RECT 190.300 116.500 190.700 116.600 ;
        RECT 192.600 116.500 193.000 116.600 ;
        RECT 190.300 116.200 193.000 116.500 ;
        RECT 189.700 115.700 192.100 115.900 ;
        RECT 194.200 115.700 194.600 119.900 ;
        RECT 189.700 115.600 194.600 115.700 ;
        RECT 191.700 115.500 194.600 115.600 ;
        RECT 191.800 115.400 194.600 115.500 ;
        RECT 195.000 115.700 195.400 119.900 ;
        RECT 197.200 118.200 197.600 119.900 ;
        RECT 196.600 117.900 197.600 118.200 ;
        RECT 199.400 117.900 199.800 119.900 ;
        RECT 201.500 117.900 202.100 119.900 ;
        RECT 196.600 117.500 197.000 117.900 ;
        RECT 199.400 117.600 199.700 117.900 ;
        RECT 198.300 117.300 200.100 117.600 ;
        RECT 201.400 117.500 201.800 117.900 ;
        RECT 198.300 117.200 198.700 117.300 ;
        RECT 199.700 117.200 200.100 117.300 ;
        RECT 196.600 116.500 197.000 116.600 ;
        RECT 198.900 116.500 199.300 116.600 ;
        RECT 196.600 116.200 199.300 116.500 ;
        RECT 199.600 116.500 200.700 116.800 ;
        RECT 199.600 115.900 199.900 116.500 ;
        RECT 200.300 116.400 200.700 116.500 ;
        RECT 201.500 116.600 202.200 117.000 ;
        RECT 201.500 116.100 201.800 116.600 ;
        RECT 197.500 115.700 199.900 115.900 ;
        RECT 195.000 115.600 199.900 115.700 ;
        RECT 200.600 115.800 201.800 116.100 ;
        RECT 195.000 115.500 197.900 115.600 ;
        RECT 195.000 115.400 197.800 115.500 ;
        RECT 186.300 114.900 186.700 115.000 ;
        RECT 186.300 114.600 188.200 114.900 ;
        RECT 188.600 114.800 189.000 115.200 ;
        RECT 191.000 115.100 191.400 115.200 ;
        RECT 198.200 115.100 198.600 115.200 ;
        RECT 191.000 114.800 193.500 115.100 ;
        RECT 187.800 114.500 188.200 114.600 ;
        RECT 188.700 114.200 189.000 114.800 ;
        RECT 193.100 114.700 193.500 114.800 ;
        RECT 196.100 114.800 198.600 115.100 ;
        RECT 196.100 114.700 196.500 114.800 ;
        RECT 197.400 114.700 197.800 114.800 ;
        RECT 192.300 114.200 192.700 114.300 ;
        RECT 196.900 114.200 197.300 114.300 ;
        RECT 200.600 114.200 200.900 115.800 ;
        RECT 203.800 115.600 204.200 119.900 ;
        RECT 202.100 115.300 204.200 115.600 ;
        RECT 202.100 115.200 202.500 115.300 ;
        RECT 202.900 114.900 203.300 115.000 ;
        RECT 201.400 114.600 203.300 114.900 ;
        RECT 201.400 114.500 201.800 114.600 ;
        RECT 188.700 114.100 194.200 114.200 ;
        RECT 195.400 114.100 200.900 114.200 ;
        RECT 188.700 113.900 200.900 114.100 ;
        RECT 188.900 113.800 189.300 113.900 ;
        RECT 185.400 113.300 187.300 113.600 ;
        RECT 183.800 111.100 184.200 113.000 ;
        RECT 185.400 111.100 185.800 113.300 ;
        RECT 186.900 113.200 187.300 113.300 ;
        RECT 191.800 112.800 192.100 113.900 ;
        RECT 193.400 113.800 196.200 113.900 ;
        RECT 190.900 112.700 191.300 112.800 ;
        RECT 187.800 112.100 188.200 112.500 ;
        RECT 189.900 112.400 191.300 112.700 ;
        RECT 191.800 112.400 192.200 112.800 ;
        RECT 189.900 112.100 190.200 112.400 ;
        RECT 192.600 112.100 193.000 112.500 ;
        RECT 187.500 111.800 188.200 112.100 ;
        RECT 187.500 111.100 188.100 111.800 ;
        RECT 189.800 111.100 190.200 112.100 ;
        RECT 192.000 111.800 193.000 112.100 ;
        RECT 192.000 111.100 192.400 111.800 ;
        RECT 194.200 111.100 194.600 113.500 ;
        RECT 195.000 111.100 195.400 113.500 ;
        RECT 197.500 112.800 197.800 113.900 ;
        RECT 200.300 113.800 200.700 113.900 ;
        RECT 203.800 113.600 204.200 115.300 ;
        RECT 202.300 113.300 204.200 113.600 ;
        RECT 202.300 113.200 202.700 113.300 ;
        RECT 196.600 112.100 197.000 112.500 ;
        RECT 197.400 112.400 197.800 112.800 ;
        RECT 198.300 112.700 198.700 112.800 ;
        RECT 198.300 112.400 199.700 112.700 ;
        RECT 199.400 112.100 199.700 112.400 ;
        RECT 201.400 112.100 201.800 112.500 ;
        RECT 196.600 111.800 197.600 112.100 ;
        RECT 197.200 111.100 197.600 111.800 ;
        RECT 199.400 111.100 199.800 112.100 ;
        RECT 201.400 111.800 202.100 112.100 ;
        RECT 201.500 111.100 202.100 111.800 ;
        RECT 203.800 111.100 204.200 113.300 ;
        RECT 0.600 107.700 1.000 109.900 ;
        RECT 2.700 109.200 3.300 109.900 ;
        RECT 2.700 108.900 3.400 109.200 ;
        RECT 5.000 108.900 5.400 109.900 ;
        RECT 7.200 109.200 7.600 109.900 ;
        RECT 7.200 108.900 8.200 109.200 ;
        RECT 3.000 108.500 3.400 108.900 ;
        RECT 5.100 108.600 5.400 108.900 ;
        RECT 5.100 108.300 6.500 108.600 ;
        RECT 6.100 108.200 6.500 108.300 ;
        RECT 7.000 108.200 7.400 108.600 ;
        RECT 7.800 108.500 8.200 108.900 ;
        RECT 2.100 107.700 2.500 107.800 ;
        RECT 0.600 107.400 2.500 107.700 ;
        RECT 0.600 105.700 1.000 107.400 ;
        RECT 4.100 107.100 4.500 107.200 ;
        RECT 6.200 107.100 6.600 107.200 ;
        RECT 7.000 107.100 7.300 108.200 ;
        RECT 9.400 107.500 9.800 109.900 ;
        RECT 10.200 107.800 10.600 108.600 ;
        RECT 8.600 107.100 9.400 107.200 ;
        RECT 3.900 106.800 9.400 107.100 ;
        RECT 3.000 106.400 3.400 106.500 ;
        RECT 1.500 106.100 3.400 106.400 ;
        RECT 1.500 106.000 1.900 106.100 ;
        RECT 2.300 105.700 2.700 105.800 ;
        RECT 0.600 105.400 2.700 105.700 ;
        RECT 0.600 101.100 1.000 105.400 ;
        RECT 3.900 105.200 4.200 106.800 ;
        RECT 7.500 106.700 7.900 106.800 ;
        RECT 7.000 106.200 7.400 106.300 ;
        RECT 8.300 106.200 8.700 106.300 ;
        RECT 6.200 105.900 8.700 106.200 ;
        RECT 6.200 105.800 6.600 105.900 ;
        RECT 7.000 105.500 9.800 105.600 ;
        RECT 6.900 105.400 9.800 105.500 ;
        RECT 3.000 104.900 4.200 105.200 ;
        RECT 4.900 105.300 9.800 105.400 ;
        RECT 4.900 105.100 7.300 105.300 ;
        RECT 3.000 104.400 3.300 104.900 ;
        RECT 2.600 104.000 3.300 104.400 ;
        RECT 4.100 104.500 4.500 104.600 ;
        RECT 4.900 104.500 5.200 105.100 ;
        RECT 4.100 104.200 5.200 104.500 ;
        RECT 5.500 104.500 8.200 104.800 ;
        RECT 5.500 104.400 5.900 104.500 ;
        RECT 7.800 104.400 8.200 104.500 ;
        RECT 4.700 103.700 5.100 103.800 ;
        RECT 6.100 103.700 6.500 103.800 ;
        RECT 3.000 103.100 3.400 103.500 ;
        RECT 4.700 103.400 6.500 103.700 ;
        RECT 5.100 103.100 5.400 103.400 ;
        RECT 7.800 103.100 8.200 103.500 ;
        RECT 2.700 101.100 3.300 103.100 ;
        RECT 5.000 101.100 5.400 103.100 ;
        RECT 7.200 102.800 8.200 103.100 ;
        RECT 7.200 101.100 7.600 102.800 ;
        RECT 9.400 101.100 9.800 105.300 ;
        RECT 11.000 101.100 11.400 109.900 ;
        RECT 11.800 108.000 12.200 109.900 ;
        RECT 13.400 108.000 13.800 109.900 ;
        RECT 11.800 107.900 13.800 108.000 ;
        RECT 14.200 107.900 14.600 109.900 ;
        RECT 15.300 108.200 15.700 109.900 ;
        RECT 19.300 109.200 19.700 109.500 ;
        RECT 19.000 108.800 19.700 109.200 ;
        RECT 15.300 107.900 16.200 108.200 ;
        RECT 19.300 108.000 19.700 108.800 ;
        RECT 21.400 108.500 21.800 109.500 ;
        RECT 11.900 107.700 13.700 107.900 ;
        RECT 12.200 107.200 12.600 107.400 ;
        RECT 14.200 107.200 14.500 107.900 ;
        RECT 11.800 106.900 12.600 107.200 ;
        RECT 11.800 106.800 12.200 106.900 ;
        RECT 13.300 106.800 14.600 107.200 ;
        RECT 12.600 105.800 13.000 106.600 ;
        RECT 13.300 105.200 13.600 106.800 ;
        RECT 15.800 106.100 16.200 107.900 ;
        RECT 18.900 107.700 19.700 108.000 ;
        RECT 16.600 107.100 17.000 107.600 ;
        RECT 18.900 107.500 19.300 107.700 ;
        RECT 18.900 107.200 19.200 107.500 ;
        RECT 21.500 107.400 21.800 108.500 ;
        RECT 22.200 107.800 22.600 108.600 ;
        RECT 17.400 107.100 17.800 107.200 ;
        RECT 16.600 106.800 17.800 107.100 ;
        RECT 18.200 106.800 19.200 107.200 ;
        RECT 19.700 107.100 21.800 107.400 ;
        RECT 19.700 106.900 20.200 107.100 ;
        RECT 12.600 104.800 13.600 105.200 ;
        RECT 14.200 105.800 16.200 106.100 ;
        RECT 16.600 106.100 17.000 106.200 ;
        RECT 17.400 106.100 17.800 106.200 ;
        RECT 18.200 106.100 18.600 106.200 ;
        RECT 16.600 105.800 18.600 106.100 ;
        RECT 14.200 105.200 14.500 105.800 ;
        RECT 14.200 105.100 14.600 105.200 ;
        RECT 13.900 104.800 14.600 105.100 ;
        RECT 13.100 101.100 13.500 104.800 ;
        RECT 13.900 104.200 14.200 104.800 ;
        RECT 15.000 104.400 15.400 105.200 ;
        RECT 13.800 103.800 14.200 104.200 ;
        RECT 15.800 101.100 16.200 105.800 ;
        RECT 18.200 105.400 18.600 105.800 ;
        RECT 18.900 104.900 19.200 106.800 ;
        RECT 19.500 106.500 20.200 106.900 ;
        RECT 19.900 105.500 20.200 106.500 ;
        RECT 20.600 105.800 21.000 106.600 ;
        RECT 21.400 105.800 21.800 106.600 ;
        RECT 23.000 106.100 23.400 109.900 ;
        RECT 23.800 108.000 24.200 109.900 ;
        RECT 25.400 108.000 25.800 109.900 ;
        RECT 23.800 107.900 25.800 108.000 ;
        RECT 26.200 107.900 26.600 109.900 ;
        RECT 23.900 107.700 25.700 107.900 ;
        RECT 24.200 107.200 24.600 107.400 ;
        RECT 26.200 107.200 26.500 107.900 ;
        RECT 27.000 107.800 27.400 108.600 ;
        RECT 23.800 106.900 24.600 107.200 ;
        RECT 23.800 106.800 24.200 106.900 ;
        RECT 25.300 106.800 26.600 107.200 ;
        RECT 24.600 106.100 25.000 106.600 ;
        RECT 23.000 105.800 25.000 106.100 ;
        RECT 25.300 106.100 25.600 106.800 ;
        RECT 26.200 106.100 26.600 106.200 ;
        RECT 25.300 105.800 26.600 106.100 ;
        RECT 19.900 105.200 21.800 105.500 ;
        RECT 18.900 104.600 19.700 104.900 ;
        RECT 19.300 101.100 19.700 104.600 ;
        RECT 21.500 103.500 21.800 105.200 ;
        RECT 21.400 101.500 21.800 103.500 ;
        RECT 23.000 101.100 23.400 105.800 ;
        RECT 25.300 105.100 25.600 105.800 ;
        RECT 26.200 105.100 26.600 105.200 ;
        RECT 25.100 104.800 25.600 105.100 ;
        RECT 25.900 104.800 26.600 105.100 ;
        RECT 25.100 101.100 25.500 104.800 ;
        RECT 25.900 104.200 26.200 104.800 ;
        RECT 25.800 103.800 26.200 104.200 ;
        RECT 27.800 101.100 28.200 109.900 ;
        RECT 30.200 107.900 30.600 109.900 ;
        RECT 30.900 108.200 31.300 108.600 ;
        RECT 29.400 106.400 29.800 107.200 ;
        RECT 28.600 106.100 29.000 106.200 ;
        RECT 30.200 106.100 30.500 107.900 ;
        RECT 31.000 107.800 31.400 108.200 ;
        RECT 31.800 107.900 32.200 109.900 ;
        RECT 32.600 108.000 33.000 109.900 ;
        RECT 34.200 108.000 34.600 109.900 ;
        RECT 32.600 107.900 34.600 108.000 ;
        RECT 31.900 107.200 32.200 107.900 ;
        RECT 32.700 107.700 34.500 107.900 ;
        RECT 35.000 107.800 35.400 108.600 ;
        RECT 33.800 107.200 34.200 107.400 ;
        RECT 31.800 106.800 33.100 107.200 ;
        RECT 33.800 106.900 34.600 107.200 ;
        RECT 34.200 106.800 34.600 106.900 ;
        RECT 31.000 106.100 31.400 106.200 ;
        RECT 28.600 105.800 29.400 106.100 ;
        RECT 30.200 105.800 31.400 106.100 ;
        RECT 31.800 106.100 32.200 106.200 ;
        RECT 32.800 106.100 33.100 106.800 ;
        RECT 31.800 105.800 33.100 106.100 ;
        RECT 33.400 105.800 33.800 106.600 ;
        RECT 29.000 105.600 29.400 105.800 ;
        RECT 31.000 105.100 31.300 105.800 ;
        RECT 31.800 105.100 32.200 105.200 ;
        RECT 32.800 105.100 33.100 105.800 ;
        RECT 28.600 104.800 30.600 105.100 ;
        RECT 28.600 101.100 29.000 104.800 ;
        RECT 30.200 101.100 30.600 104.800 ;
        RECT 31.000 104.800 32.500 105.100 ;
        RECT 32.800 104.800 33.300 105.100 ;
        RECT 31.000 101.100 31.400 104.800 ;
        RECT 32.200 104.200 32.500 104.800 ;
        RECT 32.200 103.800 32.600 104.200 ;
        RECT 32.900 101.100 33.300 104.800 ;
        RECT 35.800 101.100 36.200 109.900 ;
        RECT 36.600 108.000 37.000 109.900 ;
        RECT 38.200 108.000 38.600 109.900 ;
        RECT 36.600 107.900 38.600 108.000 ;
        RECT 39.000 107.900 39.400 109.900 ;
        RECT 39.900 108.200 40.300 108.600 ;
        RECT 36.700 107.700 38.500 107.900 ;
        RECT 37.000 107.200 37.400 107.400 ;
        RECT 39.000 107.200 39.300 107.900 ;
        RECT 39.800 107.800 40.200 108.200 ;
        RECT 40.600 107.900 41.000 109.900 ;
        RECT 36.600 106.900 37.400 107.200 ;
        RECT 36.600 106.800 37.000 106.900 ;
        RECT 38.100 106.800 39.400 107.200 ;
        RECT 36.600 106.100 37.000 106.200 ;
        RECT 37.400 106.100 37.800 106.600 ;
        RECT 36.600 105.800 37.800 106.100 ;
        RECT 38.100 106.200 38.400 106.800 ;
        RECT 38.100 105.800 38.600 106.200 ;
        RECT 39.800 106.100 40.200 106.200 ;
        RECT 40.700 106.100 41.000 107.900 ;
        RECT 44.600 107.900 45.000 109.900 ;
        RECT 45.300 108.200 45.700 108.600 ;
        RECT 47.000 108.200 47.400 109.900 ;
        RECT 41.400 106.400 41.800 107.200 ;
        RECT 43.800 106.400 44.200 107.200 ;
        RECT 42.200 106.100 42.600 106.200 ;
        RECT 39.800 105.800 41.000 106.100 ;
        RECT 41.800 105.800 42.600 106.100 ;
        RECT 43.000 106.100 43.400 106.200 ;
        RECT 44.600 106.100 44.900 107.900 ;
        RECT 45.400 107.800 45.800 108.200 ;
        RECT 46.900 107.900 47.400 108.200 ;
        RECT 46.900 107.200 47.200 107.900 ;
        RECT 48.600 107.600 49.000 109.900 ;
        RECT 47.700 107.300 49.000 107.600 ;
        RECT 51.000 107.600 51.400 109.900 ;
        RECT 52.600 108.200 53.000 109.900 ;
        RECT 55.000 108.200 55.400 109.900 ;
        RECT 52.600 107.900 53.100 108.200 ;
        RECT 51.000 107.300 52.300 107.600 ;
        RECT 46.200 107.100 46.600 107.200 ;
        RECT 46.900 107.100 47.400 107.200 ;
        RECT 46.200 106.800 47.400 107.100 ;
        RECT 45.400 106.100 45.800 106.200 ;
        RECT 43.000 105.800 43.800 106.100 ;
        RECT 44.600 105.800 45.800 106.100 ;
        RECT 38.100 105.100 38.400 105.800 ;
        RECT 39.000 105.100 39.400 105.200 ;
        RECT 39.900 105.100 40.200 105.800 ;
        RECT 41.800 105.600 42.200 105.800 ;
        RECT 43.400 105.600 43.800 105.800 ;
        RECT 45.400 105.100 45.700 105.800 ;
        RECT 46.900 105.100 47.200 106.800 ;
        RECT 47.700 106.500 48.000 107.300 ;
        RECT 47.500 106.100 48.000 106.500 ;
        RECT 47.700 105.100 48.000 106.100 ;
        RECT 48.500 106.200 48.900 106.600 ;
        RECT 51.100 106.200 51.500 106.600 ;
        RECT 48.500 106.100 49.000 106.200 ;
        RECT 51.000 106.100 51.500 106.200 ;
        RECT 48.500 105.800 51.500 106.100 ;
        RECT 52.000 106.500 52.300 107.300 ;
        RECT 52.800 107.200 53.100 107.900 ;
        RECT 52.600 106.800 53.100 107.200 ;
        RECT 52.000 106.100 52.500 106.500 ;
        RECT 52.000 105.100 52.300 106.100 ;
        RECT 52.800 105.100 53.100 106.800 ;
        RECT 37.900 104.800 38.400 105.100 ;
        RECT 38.700 104.800 40.200 105.100 ;
        RECT 37.900 101.100 38.300 104.800 ;
        RECT 38.700 104.200 39.000 104.800 ;
        RECT 38.600 103.800 39.000 104.200 ;
        RECT 39.800 101.100 40.200 104.800 ;
        RECT 40.600 104.800 42.600 105.100 ;
        RECT 40.600 101.100 41.000 104.800 ;
        RECT 42.200 101.100 42.600 104.800 ;
        RECT 43.000 104.800 45.000 105.100 ;
        RECT 43.000 101.100 43.400 104.800 ;
        RECT 44.600 101.100 45.000 104.800 ;
        RECT 45.400 101.100 45.800 105.100 ;
        RECT 46.900 104.600 47.400 105.100 ;
        RECT 47.700 104.800 49.000 105.100 ;
        RECT 47.000 101.100 47.400 104.600 ;
        RECT 48.600 101.100 49.000 104.800 ;
        RECT 51.000 104.800 52.300 105.100 ;
        RECT 51.000 101.100 51.400 104.800 ;
        RECT 52.600 104.600 53.100 105.100 ;
        RECT 54.900 107.900 55.400 108.200 ;
        RECT 54.900 107.200 55.200 107.900 ;
        RECT 56.600 107.600 57.000 109.900 ;
        RECT 57.400 109.600 59.400 109.900 ;
        RECT 57.400 107.900 57.800 109.600 ;
        RECT 58.200 107.900 58.600 109.300 ;
        RECT 59.000 108.000 59.400 109.600 ;
        RECT 60.600 108.000 61.000 109.900 ;
        RECT 62.200 108.200 62.600 109.900 ;
        RECT 59.000 107.900 61.000 108.000 ;
        RECT 62.100 107.900 62.600 108.200 ;
        RECT 55.700 107.300 57.000 107.600 ;
        RECT 54.900 106.800 55.400 107.200 ;
        RECT 54.900 105.100 55.200 106.800 ;
        RECT 55.700 106.500 56.000 107.300 ;
        RECT 58.200 107.200 58.500 107.900 ;
        RECT 59.100 107.700 60.900 107.900 ;
        RECT 60.200 107.200 60.600 107.400 ;
        RECT 62.100 107.200 62.400 107.900 ;
        RECT 63.800 107.600 64.200 109.900 ;
        RECT 64.600 107.800 65.000 108.600 ;
        RECT 62.900 107.300 64.200 107.600 ;
        RECT 55.500 106.100 56.000 106.500 ;
        RECT 55.700 105.100 56.000 106.100 ;
        RECT 56.500 106.200 56.900 106.600 ;
        RECT 57.400 106.400 57.800 107.200 ;
        RECT 58.200 106.900 59.400 107.200 ;
        RECT 60.200 106.900 61.000 107.200 ;
        RECT 59.000 106.800 59.400 106.900 ;
        RECT 60.600 106.800 61.000 106.900 ;
        RECT 61.400 107.100 61.800 107.200 ;
        RECT 62.100 107.100 62.600 107.200 ;
        RECT 61.400 106.800 62.600 107.100 ;
        RECT 56.500 105.800 57.000 106.200 ;
        RECT 58.200 105.800 58.600 106.600 ;
        RECT 59.100 105.100 59.400 106.800 ;
        RECT 59.800 105.800 60.200 106.600 ;
        RECT 62.100 105.100 62.400 106.800 ;
        RECT 62.900 106.500 63.200 107.300 ;
        RECT 62.700 106.100 63.200 106.500 ;
        RECT 62.900 105.100 63.200 106.100 ;
        RECT 63.700 106.200 64.100 106.600 ;
        RECT 63.700 105.800 64.200 106.200 ;
        RECT 54.900 104.600 55.400 105.100 ;
        RECT 55.700 104.800 57.000 105.100 ;
        RECT 52.600 101.100 53.000 104.600 ;
        RECT 55.000 101.100 55.400 104.600 ;
        RECT 56.600 101.100 57.000 104.800 ;
        RECT 58.700 101.100 59.700 105.100 ;
        RECT 62.100 104.600 62.600 105.100 ;
        RECT 62.900 104.800 64.200 105.100 ;
        RECT 62.200 101.100 62.600 104.600 ;
        RECT 63.800 101.100 64.200 104.800 ;
        RECT 65.400 101.100 65.800 109.900 ;
        RECT 66.300 108.200 66.700 108.600 ;
        RECT 66.200 107.800 66.600 108.200 ;
        RECT 67.000 107.900 67.400 109.900 ;
        RECT 69.400 108.000 69.800 109.900 ;
        RECT 71.000 109.600 73.000 109.900 ;
        RECT 71.000 108.000 71.400 109.600 ;
        RECT 69.400 107.900 71.400 108.000 ;
        RECT 71.800 107.900 72.200 109.300 ;
        RECT 72.600 107.900 73.000 109.600 ;
        RECT 74.200 108.900 74.600 109.900 ;
        RECT 66.200 106.100 66.600 106.200 ;
        RECT 67.100 106.100 67.400 107.900 ;
        RECT 69.500 107.700 71.300 107.900 ;
        RECT 69.800 107.200 70.200 107.400 ;
        RECT 71.900 107.200 72.200 107.900 ;
        RECT 73.400 107.800 73.800 108.600 ;
        RECT 74.300 107.200 74.600 108.900 ;
        RECT 75.800 107.500 76.200 109.900 ;
        RECT 78.000 109.200 78.400 109.900 ;
        RECT 77.400 108.900 78.400 109.200 ;
        RECT 80.200 108.900 80.600 109.900 ;
        RECT 82.300 109.200 82.900 109.900 ;
        RECT 82.200 108.900 82.900 109.200 ;
        RECT 77.400 108.500 77.800 108.900 ;
        RECT 80.200 108.600 80.500 108.900 ;
        RECT 78.200 107.800 78.600 108.600 ;
        RECT 79.100 108.300 80.500 108.600 ;
        RECT 82.200 108.500 82.600 108.900 ;
        RECT 79.100 108.200 79.500 108.300 ;
        RECT 67.800 106.400 68.200 107.200 ;
        RECT 69.400 106.900 70.200 107.200 ;
        RECT 71.000 106.900 72.200 107.200 ;
        RECT 69.400 106.800 69.800 106.900 ;
        RECT 71.000 106.800 71.400 106.900 ;
        RECT 68.600 106.100 69.000 106.200 ;
        RECT 66.200 105.800 67.400 106.100 ;
        RECT 68.200 105.800 69.000 106.100 ;
        RECT 70.200 105.800 70.600 106.600 ;
        RECT 66.300 105.100 66.600 105.800 ;
        RECT 68.200 105.600 68.600 105.800 ;
        RECT 71.000 105.100 71.300 106.800 ;
        RECT 71.800 105.800 72.200 106.600 ;
        RECT 72.600 106.400 73.000 107.200 ;
        RECT 74.200 106.800 74.600 107.200 ;
        RECT 76.200 107.100 77.000 107.200 ;
        RECT 78.300 107.100 78.600 107.800 ;
        RECT 83.100 107.700 83.500 107.800 ;
        RECT 84.600 107.700 85.000 109.900 ;
        RECT 85.700 108.200 86.100 109.900 ;
        RECT 88.600 108.900 89.000 109.900 ;
        RECT 85.700 107.900 86.600 108.200 ;
        RECT 83.100 107.400 85.000 107.700 ;
        RECT 81.100 107.100 81.500 107.200 ;
        RECT 76.200 106.800 81.700 107.100 ;
        RECT 74.300 105.100 74.600 106.800 ;
        RECT 77.700 106.700 78.100 106.800 ;
        RECT 76.900 106.200 77.300 106.300 ;
        RECT 75.000 105.400 75.400 106.200 ;
        RECT 76.900 106.100 79.400 106.200 ;
        RECT 79.800 106.100 80.200 106.200 ;
        RECT 76.900 105.900 80.200 106.100 ;
        RECT 79.000 105.800 80.200 105.900 ;
        RECT 75.800 105.500 78.600 105.600 ;
        RECT 75.800 105.400 78.700 105.500 ;
        RECT 75.800 105.300 80.700 105.400 ;
        RECT 66.200 101.100 66.600 105.100 ;
        RECT 67.000 104.800 69.000 105.100 ;
        RECT 67.000 101.100 67.400 104.800 ;
        RECT 68.600 101.100 69.000 104.800 ;
        RECT 70.700 101.100 71.700 105.100 ;
        RECT 74.200 104.700 75.100 105.100 ;
        RECT 74.700 102.200 75.100 104.700 ;
        RECT 74.200 101.800 75.100 102.200 ;
        RECT 74.700 101.100 75.100 101.800 ;
        RECT 75.800 101.100 76.200 105.300 ;
        RECT 78.300 105.100 80.700 105.300 ;
        RECT 77.400 104.500 80.100 104.800 ;
        RECT 77.400 104.400 77.800 104.500 ;
        RECT 79.700 104.400 80.100 104.500 ;
        RECT 80.400 104.500 80.700 105.100 ;
        RECT 81.400 105.200 81.700 106.800 ;
        RECT 82.200 106.400 82.600 106.500 ;
        RECT 82.200 106.100 84.100 106.400 ;
        RECT 83.700 106.000 84.100 106.100 ;
        RECT 82.900 105.700 83.300 105.800 ;
        RECT 84.600 105.700 85.000 107.400 ;
        RECT 85.400 106.800 85.800 107.200 ;
        RECT 85.400 106.100 85.700 106.800 ;
        RECT 86.200 106.100 86.600 107.900 ;
        RECT 87.000 106.800 87.400 107.600 ;
        RECT 88.600 107.200 88.900 108.900 ;
        RECT 89.400 107.800 89.800 108.600 ;
        RECT 90.200 107.900 90.600 109.900 ;
        RECT 91.000 108.000 91.400 109.900 ;
        RECT 92.600 108.000 93.000 109.900 ;
        RECT 94.200 108.200 94.600 109.900 ;
        RECT 91.000 107.900 93.000 108.000 ;
        RECT 90.300 107.200 90.600 107.900 ;
        RECT 91.100 107.700 92.900 107.900 ;
        RECT 94.100 107.800 94.600 108.200 ;
        RECT 92.200 107.200 92.600 107.400 ;
        RECT 94.100 107.200 94.400 107.800 ;
        RECT 95.800 107.600 96.200 109.900 ;
        RECT 94.900 107.300 96.200 107.600 ;
        RECT 88.600 106.800 89.000 107.200 ;
        RECT 90.200 107.100 91.500 107.200 ;
        RECT 89.400 106.800 91.500 107.100 ;
        RECT 92.200 106.900 93.000 107.200 ;
        RECT 92.600 106.800 93.000 106.900 ;
        RECT 94.100 106.800 94.600 107.200 ;
        RECT 85.400 105.800 86.600 106.100 ;
        RECT 82.900 105.400 85.000 105.700 ;
        RECT 81.400 104.900 82.600 105.200 ;
        RECT 81.100 104.500 81.500 104.600 ;
        RECT 80.400 104.200 81.500 104.500 ;
        RECT 82.300 104.400 82.600 104.900 ;
        RECT 82.300 104.000 83.000 104.400 ;
        RECT 79.100 103.700 79.500 103.800 ;
        RECT 80.500 103.700 80.900 103.800 ;
        RECT 77.400 103.100 77.800 103.500 ;
        RECT 79.100 103.400 80.900 103.700 ;
        RECT 80.200 103.100 80.500 103.400 ;
        RECT 82.200 103.100 82.600 103.500 ;
        RECT 77.400 102.800 78.400 103.100 ;
        RECT 78.000 101.100 78.400 102.800 ;
        RECT 80.200 101.100 80.600 103.100 ;
        RECT 82.300 101.100 82.900 103.100 ;
        RECT 84.600 101.100 85.000 105.400 ;
        RECT 85.400 104.400 85.800 105.200 ;
        RECT 86.200 101.100 86.600 105.800 ;
        RECT 87.800 105.400 88.200 106.200 ;
        RECT 88.600 105.100 88.900 106.800 ;
        RECT 89.400 106.200 89.700 106.800 ;
        RECT 89.400 105.800 89.800 106.200 ;
        RECT 90.200 105.100 90.600 105.200 ;
        RECT 91.200 105.100 91.500 106.800 ;
        RECT 91.800 105.800 92.200 106.600 ;
        RECT 94.100 105.100 94.400 106.800 ;
        RECT 94.900 106.500 95.200 107.300 ;
        RECT 94.700 106.100 95.200 106.500 ;
        RECT 94.900 105.100 95.200 106.100 ;
        RECT 95.700 106.200 96.100 106.600 ;
        RECT 95.700 105.800 96.200 106.200 ;
        RECT 88.100 104.700 89.000 105.100 ;
        RECT 90.200 104.800 90.900 105.100 ;
        RECT 91.200 104.800 91.700 105.100 ;
        RECT 88.100 102.200 88.500 104.700 ;
        RECT 90.600 104.200 90.900 104.800 ;
        RECT 90.600 103.800 91.000 104.200 ;
        RECT 88.100 101.800 89.000 102.200 ;
        RECT 88.100 101.100 88.500 101.800 ;
        RECT 91.300 101.100 91.700 104.800 ;
        RECT 94.100 104.600 94.600 105.100 ;
        RECT 94.900 104.800 96.200 105.100 ;
        RECT 94.200 101.100 94.600 104.600 ;
        RECT 95.800 101.100 96.200 104.800 ;
        RECT 96.600 101.100 97.000 109.900 ;
        RECT 97.400 107.800 97.800 108.600 ;
        RECT 99.500 108.200 99.900 109.900 ;
        RECT 99.000 107.900 99.900 108.200 ;
        RECT 102.200 107.900 102.600 109.900 ;
        RECT 103.000 108.000 103.400 109.900 ;
        RECT 104.600 108.000 105.000 109.900 ;
        RECT 103.000 107.900 105.000 108.000 ;
        RECT 98.200 106.800 98.600 107.600 ;
        RECT 99.000 106.100 99.400 107.900 ;
        RECT 102.300 107.200 102.600 107.900 ;
        RECT 103.100 107.700 104.900 107.900 ;
        RECT 105.400 107.700 105.800 109.900 ;
        RECT 107.500 109.200 108.100 109.900 ;
        RECT 107.500 108.900 108.200 109.200 ;
        RECT 109.800 108.900 110.200 109.900 ;
        RECT 112.000 109.200 112.400 109.900 ;
        RECT 112.000 108.900 113.000 109.200 ;
        RECT 107.800 108.500 108.200 108.900 ;
        RECT 109.900 108.600 110.200 108.900 ;
        RECT 109.900 108.300 111.300 108.600 ;
        RECT 110.900 108.200 111.300 108.300 ;
        RECT 111.800 108.200 112.200 108.600 ;
        RECT 112.600 108.500 113.000 108.900 ;
        RECT 106.900 107.700 107.300 107.800 ;
        RECT 105.400 107.400 107.300 107.700 ;
        RECT 104.200 107.200 104.600 107.400 ;
        RECT 102.200 106.800 103.500 107.200 ;
        RECT 104.200 106.900 105.000 107.200 ;
        RECT 104.600 106.800 105.000 106.900 ;
        RECT 103.200 106.200 103.500 106.800 ;
        RECT 99.000 105.800 102.500 106.100 ;
        RECT 103.000 105.800 103.500 106.200 ;
        RECT 103.800 105.800 104.200 106.600 ;
        RECT 99.000 101.100 99.400 105.800 ;
        RECT 102.200 105.200 102.500 105.800 ;
        RECT 99.800 104.400 100.200 105.200 ;
        RECT 102.200 105.100 102.600 105.200 ;
        RECT 103.200 105.100 103.500 105.800 ;
        RECT 105.400 105.700 105.800 107.400 ;
        RECT 108.900 107.100 109.300 107.200 ;
        RECT 111.800 107.100 112.100 108.200 ;
        RECT 114.200 107.500 114.600 109.900 ;
        RECT 115.000 107.600 115.400 109.900 ;
        RECT 116.600 108.200 117.000 109.900 ;
        RECT 116.600 107.900 117.100 108.200 ;
        RECT 115.000 107.300 116.300 107.600 ;
        RECT 113.400 107.100 114.200 107.200 ;
        RECT 108.700 106.800 114.200 107.100 ;
        RECT 107.800 106.400 108.200 106.500 ;
        RECT 106.300 106.100 108.200 106.400 ;
        RECT 106.300 106.000 106.700 106.100 ;
        RECT 107.100 105.700 107.500 105.800 ;
        RECT 105.400 105.400 107.500 105.700 ;
        RECT 102.200 104.800 102.900 105.100 ;
        RECT 103.200 104.800 103.700 105.100 ;
        RECT 102.600 104.200 102.900 104.800 ;
        RECT 102.600 103.800 103.000 104.200 ;
        RECT 103.300 101.100 103.700 104.800 ;
        RECT 105.400 101.100 105.800 105.400 ;
        RECT 108.700 105.200 109.000 106.800 ;
        RECT 112.300 106.700 112.700 106.800 ;
        RECT 113.100 106.200 113.500 106.300 ;
        RECT 115.100 106.200 115.500 106.600 ;
        RECT 111.000 105.900 113.500 106.200 ;
        RECT 111.000 105.800 111.400 105.900 ;
        RECT 115.000 105.800 115.500 106.200 ;
        RECT 116.000 106.500 116.300 107.300 ;
        RECT 116.800 107.200 117.100 107.900 ;
        RECT 118.200 107.500 118.600 109.900 ;
        RECT 120.400 109.200 120.800 109.900 ;
        RECT 119.800 108.900 120.800 109.200 ;
        RECT 122.600 108.900 123.000 109.900 ;
        RECT 124.700 109.200 125.300 109.900 ;
        RECT 124.600 108.900 125.300 109.200 ;
        RECT 119.800 108.500 120.200 108.900 ;
        RECT 122.600 108.600 122.900 108.900 ;
        RECT 120.600 107.800 121.000 108.600 ;
        RECT 121.500 108.300 122.900 108.600 ;
        RECT 124.600 108.500 125.000 108.900 ;
        RECT 121.500 108.200 121.900 108.300 ;
        RECT 127.000 108.100 127.400 109.900 ;
        RECT 128.600 108.900 129.000 109.900 ;
        RECT 127.800 108.100 128.200 108.600 ;
        RECT 128.700 108.100 129.000 108.900 ;
        RECT 130.300 108.200 130.700 108.600 ;
        RECT 130.200 108.100 130.600 108.200 ;
        RECT 127.000 107.800 128.200 108.100 ;
        RECT 128.600 107.800 130.600 108.100 ;
        RECT 131.000 107.900 131.400 109.900 ;
        RECT 116.600 106.800 117.100 107.200 ;
        RECT 118.600 107.100 119.400 107.200 ;
        RECT 120.700 107.100 121.000 107.800 ;
        RECT 125.500 107.700 125.900 107.800 ;
        RECT 127.000 107.700 127.400 107.800 ;
        RECT 125.500 107.400 127.400 107.700 ;
        RECT 123.500 107.100 123.900 107.200 ;
        RECT 118.600 106.800 124.100 107.100 ;
        RECT 116.000 106.100 116.500 106.500 ;
        RECT 111.800 105.500 114.600 105.600 ;
        RECT 111.700 105.400 114.600 105.500 ;
        RECT 107.800 104.900 109.000 105.200 ;
        RECT 109.700 105.300 114.600 105.400 ;
        RECT 109.700 105.100 112.100 105.300 ;
        RECT 107.800 104.400 108.100 104.900 ;
        RECT 107.400 104.000 108.100 104.400 ;
        RECT 108.900 104.500 109.300 104.600 ;
        RECT 109.700 104.500 110.000 105.100 ;
        RECT 108.900 104.200 110.000 104.500 ;
        RECT 110.300 104.500 113.000 104.800 ;
        RECT 110.300 104.400 110.700 104.500 ;
        RECT 112.600 104.400 113.000 104.500 ;
        RECT 109.500 103.700 109.900 103.800 ;
        RECT 110.900 103.700 111.300 103.800 ;
        RECT 107.800 103.100 108.200 103.500 ;
        RECT 109.500 103.400 111.300 103.700 ;
        RECT 109.900 103.100 110.200 103.400 ;
        RECT 112.600 103.100 113.000 103.500 ;
        RECT 107.500 101.100 108.100 103.100 ;
        RECT 109.800 101.100 110.200 103.100 ;
        RECT 112.000 102.800 113.000 103.100 ;
        RECT 112.000 101.100 112.400 102.800 ;
        RECT 114.200 101.100 114.600 105.300 ;
        RECT 116.000 105.100 116.300 106.100 ;
        RECT 116.800 105.100 117.100 106.800 ;
        RECT 120.100 106.700 120.500 106.800 ;
        RECT 119.300 106.200 119.700 106.300 ;
        RECT 119.300 105.900 121.800 106.200 ;
        RECT 121.400 105.800 121.800 105.900 ;
        RECT 115.000 104.800 116.300 105.100 ;
        RECT 115.000 101.100 115.400 104.800 ;
        RECT 116.600 104.600 117.100 105.100 ;
        RECT 118.200 105.500 121.000 105.600 ;
        RECT 118.200 105.400 121.100 105.500 ;
        RECT 118.200 105.300 123.100 105.400 ;
        RECT 116.600 101.100 117.000 104.600 ;
        RECT 118.200 101.100 118.600 105.300 ;
        RECT 120.700 105.100 123.100 105.300 ;
        RECT 119.800 104.500 122.500 104.800 ;
        RECT 119.800 104.400 120.200 104.500 ;
        RECT 122.100 104.400 122.500 104.500 ;
        RECT 122.800 104.500 123.100 105.100 ;
        RECT 123.800 105.200 124.100 106.800 ;
        RECT 124.600 106.400 125.000 106.500 ;
        RECT 124.600 106.100 126.500 106.400 ;
        RECT 126.100 106.000 126.500 106.100 ;
        RECT 125.300 105.700 125.700 105.800 ;
        RECT 127.000 105.700 127.400 107.400 ;
        RECT 128.700 107.200 129.000 107.800 ;
        RECT 128.600 106.800 129.000 107.200 ;
        RECT 125.300 105.400 127.400 105.700 ;
        RECT 123.800 104.900 125.000 105.200 ;
        RECT 123.500 104.500 123.900 104.600 ;
        RECT 122.800 104.200 123.900 104.500 ;
        RECT 124.700 104.400 125.000 104.900 ;
        RECT 124.700 104.000 125.400 104.400 ;
        RECT 121.500 103.700 121.900 103.800 ;
        RECT 122.900 103.700 123.300 103.800 ;
        RECT 119.800 103.100 120.200 103.500 ;
        RECT 121.500 103.400 123.300 103.700 ;
        RECT 122.600 103.100 122.900 103.400 ;
        RECT 124.600 103.100 125.000 103.500 ;
        RECT 119.800 102.800 120.800 103.100 ;
        RECT 120.400 101.100 120.800 102.800 ;
        RECT 122.600 101.100 123.000 103.100 ;
        RECT 124.700 101.100 125.300 103.100 ;
        RECT 127.000 101.100 127.400 105.400 ;
        RECT 128.700 105.100 129.000 106.800 ;
        RECT 129.400 105.400 129.800 106.200 ;
        RECT 130.200 106.100 130.600 106.200 ;
        RECT 131.100 106.100 131.400 107.900 ;
        RECT 133.400 108.500 133.800 109.500 ;
        RECT 133.400 107.400 133.700 108.500 ;
        RECT 135.500 108.000 135.900 109.500 ;
        RECT 135.500 107.700 136.300 108.000 ;
        RECT 135.900 107.500 136.300 107.700 ;
        RECT 131.800 106.400 132.200 107.200 ;
        RECT 133.400 107.100 135.500 107.400 ;
        RECT 135.000 106.900 135.500 107.100 ;
        RECT 136.000 107.200 136.300 107.500 ;
        RECT 136.000 107.100 137.000 107.200 ;
        RECT 137.400 107.100 137.800 107.200 ;
        RECT 132.600 106.100 133.000 106.200 ;
        RECT 130.200 105.800 131.400 106.100 ;
        RECT 132.200 105.800 133.000 106.100 ;
        RECT 133.400 105.800 133.800 106.600 ;
        RECT 134.200 105.800 134.600 106.600 ;
        RECT 135.000 106.500 135.700 106.900 ;
        RECT 136.000 106.800 137.800 107.100 ;
        RECT 130.300 105.100 130.600 105.800 ;
        RECT 132.200 105.600 132.600 105.800 ;
        RECT 135.000 105.500 135.300 106.500 ;
        RECT 133.400 105.200 135.300 105.500 ;
        RECT 128.600 104.700 129.500 105.100 ;
        RECT 129.100 101.100 129.500 104.700 ;
        RECT 130.200 101.100 130.600 105.100 ;
        RECT 131.000 104.800 133.000 105.100 ;
        RECT 131.000 101.100 131.400 104.800 ;
        RECT 132.600 101.100 133.000 104.800 ;
        RECT 133.400 103.500 133.700 105.200 ;
        RECT 136.000 104.900 136.300 106.800 ;
        RECT 136.600 105.400 137.000 106.200 ;
        RECT 135.500 104.600 136.300 104.900 ;
        RECT 133.400 101.500 133.800 103.500 ;
        RECT 135.500 101.100 135.900 104.600 ;
        RECT 138.200 101.100 138.600 109.900 ;
        RECT 139.000 108.100 139.400 108.600 ;
        RECT 139.800 108.100 140.200 109.900 ;
        RECT 141.900 109.200 142.500 109.900 ;
        RECT 141.900 108.900 142.600 109.200 ;
        RECT 144.200 108.900 144.600 109.900 ;
        RECT 146.400 109.200 146.800 109.900 ;
        RECT 146.400 108.900 147.400 109.200 ;
        RECT 142.200 108.500 142.600 108.900 ;
        RECT 144.300 108.600 144.600 108.900 ;
        RECT 144.300 108.300 145.700 108.600 ;
        RECT 145.300 108.200 145.700 108.300 ;
        RECT 146.200 108.200 146.600 108.600 ;
        RECT 147.000 108.500 147.400 108.900 ;
        RECT 139.000 107.800 140.200 108.100 ;
        RECT 139.800 107.700 140.200 107.800 ;
        RECT 141.300 107.700 141.700 107.800 ;
        RECT 139.800 107.400 141.700 107.700 ;
        RECT 139.800 105.700 140.200 107.400 ;
        RECT 143.300 107.100 143.700 107.200 ;
        RECT 146.200 107.100 146.500 108.200 ;
        RECT 148.600 107.500 149.000 109.900 ;
        RECT 151.000 107.500 151.400 109.900 ;
        RECT 153.200 109.200 153.600 109.900 ;
        RECT 152.600 108.900 153.600 109.200 ;
        RECT 155.400 108.900 155.800 109.900 ;
        RECT 157.500 109.200 158.100 109.900 ;
        RECT 157.400 108.900 158.100 109.200 ;
        RECT 152.600 108.500 153.000 108.900 ;
        RECT 155.400 108.600 155.700 108.900 ;
        RECT 153.400 108.200 153.800 108.600 ;
        RECT 154.300 108.300 155.700 108.600 ;
        RECT 157.400 108.500 157.800 108.900 ;
        RECT 154.300 108.200 154.700 108.300 ;
        RECT 147.800 107.100 148.600 107.200 ;
        RECT 151.400 107.100 152.200 107.200 ;
        RECT 153.500 107.100 153.800 108.200 ;
        RECT 158.300 107.700 158.700 107.800 ;
        RECT 159.800 107.700 160.200 109.900 ;
        RECT 158.300 107.400 160.200 107.700 ;
        RECT 156.300 107.100 156.700 107.200 ;
        RECT 143.100 106.800 156.900 107.100 ;
        RECT 142.200 106.400 142.600 106.500 ;
        RECT 140.700 106.100 142.600 106.400 ;
        RECT 140.700 106.000 141.100 106.100 ;
        RECT 141.500 105.700 141.900 105.800 ;
        RECT 139.800 105.400 141.900 105.700 ;
        RECT 139.800 101.100 140.200 105.400 ;
        RECT 143.100 105.200 143.400 106.800 ;
        RECT 146.700 106.700 147.100 106.800 ;
        RECT 152.900 106.700 153.300 106.800 ;
        RECT 147.500 106.200 147.900 106.300 ;
        RECT 145.400 105.900 147.900 106.200 ;
        RECT 152.100 106.200 152.500 106.300 ;
        RECT 152.100 106.100 154.600 106.200 ;
        RECT 155.800 106.100 156.200 106.200 ;
        RECT 152.100 105.900 156.200 106.100 ;
        RECT 145.400 105.800 145.800 105.900 ;
        RECT 154.200 105.800 156.200 105.900 ;
        RECT 146.200 105.500 149.000 105.600 ;
        RECT 146.100 105.400 149.000 105.500 ;
        RECT 142.200 104.900 143.400 105.200 ;
        RECT 144.100 105.300 149.000 105.400 ;
        RECT 144.100 105.100 146.500 105.300 ;
        RECT 142.200 104.400 142.500 104.900 ;
        RECT 141.800 104.000 142.500 104.400 ;
        RECT 143.300 104.500 143.700 104.600 ;
        RECT 144.100 104.500 144.400 105.100 ;
        RECT 143.300 104.200 144.400 104.500 ;
        RECT 144.700 104.500 147.400 104.800 ;
        RECT 144.700 104.400 145.100 104.500 ;
        RECT 147.000 104.400 147.400 104.500 ;
        RECT 143.900 103.700 144.300 103.800 ;
        RECT 145.300 103.700 145.700 103.800 ;
        RECT 142.200 103.100 142.600 103.500 ;
        RECT 143.900 103.400 145.700 103.700 ;
        RECT 144.300 103.100 144.600 103.400 ;
        RECT 147.000 103.100 147.400 103.500 ;
        RECT 141.900 101.100 142.500 103.100 ;
        RECT 144.200 101.100 144.600 103.100 ;
        RECT 146.400 102.800 147.400 103.100 ;
        RECT 146.400 101.100 146.800 102.800 ;
        RECT 148.600 101.100 149.000 105.300 ;
        RECT 151.000 105.500 153.800 105.600 ;
        RECT 151.000 105.400 153.900 105.500 ;
        RECT 151.000 105.300 155.900 105.400 ;
        RECT 151.000 101.100 151.400 105.300 ;
        RECT 153.500 105.100 155.900 105.300 ;
        RECT 152.600 104.500 155.300 104.800 ;
        RECT 152.600 104.400 153.000 104.500 ;
        RECT 154.900 104.400 155.300 104.500 ;
        RECT 155.600 104.500 155.900 105.100 ;
        RECT 156.600 105.200 156.900 106.800 ;
        RECT 157.400 106.400 157.800 106.500 ;
        RECT 157.400 106.100 159.300 106.400 ;
        RECT 158.900 106.000 159.300 106.100 ;
        RECT 158.100 105.700 158.500 105.800 ;
        RECT 159.800 105.700 160.200 107.400 ;
        RECT 162.200 107.900 162.600 109.900 ;
        RECT 164.600 108.900 165.000 109.900 ;
        RECT 162.900 108.200 163.300 108.600 ;
        RECT 163.000 108.100 163.400 108.200 ;
        RECT 164.600 108.100 164.900 108.900 ;
        RECT 161.400 106.400 161.800 107.200 ;
        RECT 160.600 106.100 161.000 106.200 ;
        RECT 162.200 106.100 162.500 107.900 ;
        RECT 163.000 107.800 164.900 108.100 ;
        RECT 164.600 107.200 164.900 107.800 ;
        RECT 165.400 107.800 165.800 108.600 ;
        RECT 167.800 107.800 168.200 109.900 ;
        RECT 168.500 108.200 168.900 108.600 ;
        RECT 168.600 107.800 169.000 108.200 ;
        RECT 164.600 106.800 165.000 107.200 ;
        RECT 165.400 107.100 165.700 107.800 ;
        RECT 167.000 107.100 167.400 107.200 ;
        RECT 165.400 106.800 167.400 107.100 ;
        RECT 163.000 106.100 163.400 106.200 ;
        RECT 160.600 105.800 161.400 106.100 ;
        RECT 162.200 105.800 163.400 106.100 ;
        RECT 158.100 105.400 160.200 105.700 ;
        RECT 161.000 105.600 161.400 105.800 ;
        RECT 156.600 104.900 157.800 105.200 ;
        RECT 156.300 104.500 156.700 104.600 ;
        RECT 155.600 104.200 156.700 104.500 ;
        RECT 157.500 104.400 157.800 104.900 ;
        RECT 157.500 104.000 158.200 104.400 ;
        RECT 154.300 103.700 154.700 103.800 ;
        RECT 155.700 103.700 156.100 103.800 ;
        RECT 152.600 103.100 153.000 103.500 ;
        RECT 154.300 103.400 156.100 103.700 ;
        RECT 155.400 103.100 155.700 103.400 ;
        RECT 157.400 103.100 157.800 103.500 ;
        RECT 152.600 102.800 153.600 103.100 ;
        RECT 153.200 101.100 153.600 102.800 ;
        RECT 155.400 101.100 155.800 103.100 ;
        RECT 157.500 101.100 158.100 103.100 ;
        RECT 159.800 101.100 160.200 105.400 ;
        RECT 163.000 105.100 163.300 105.800 ;
        RECT 163.800 105.400 164.200 106.200 ;
        RECT 164.600 105.100 164.900 106.800 ;
        RECT 167.000 106.400 167.400 106.800 ;
        RECT 166.200 106.100 166.600 106.200 ;
        RECT 167.800 106.100 168.100 107.800 ;
        RECT 169.400 107.600 169.800 109.900 ;
        RECT 171.000 108.200 171.400 109.900 ;
        RECT 171.000 107.800 171.500 108.200 ;
        RECT 172.600 107.900 173.000 109.900 ;
        RECT 173.400 108.000 173.800 109.900 ;
        RECT 175.000 108.000 175.400 109.900 ;
        RECT 173.400 107.900 175.400 108.000 ;
        RECT 169.400 107.300 170.700 107.600 ;
        RECT 169.500 106.200 169.900 106.600 ;
        RECT 168.600 106.100 169.000 106.200 ;
        RECT 166.200 105.800 167.000 106.100 ;
        RECT 167.800 105.800 169.000 106.100 ;
        RECT 169.400 105.800 169.900 106.200 ;
        RECT 170.400 106.500 170.700 107.300 ;
        RECT 171.200 107.200 171.500 107.800 ;
        RECT 172.700 107.200 173.000 107.900 ;
        RECT 173.500 107.700 175.300 107.900 ;
        RECT 174.600 107.200 175.000 107.400 ;
        RECT 171.000 106.800 171.500 107.200 ;
        RECT 172.600 106.800 173.900 107.200 ;
        RECT 174.600 106.900 175.400 107.200 ;
        RECT 175.000 106.800 175.400 106.900 ;
        RECT 170.400 106.100 170.900 106.500 ;
        RECT 166.600 105.600 167.000 105.800 ;
        RECT 168.600 105.100 168.900 105.800 ;
        RECT 170.400 105.100 170.700 106.100 ;
        RECT 171.200 105.100 171.500 106.800 ;
        RECT 160.600 104.800 162.600 105.100 ;
        RECT 160.600 101.100 161.000 104.800 ;
        RECT 162.200 101.100 162.600 104.800 ;
        RECT 163.000 101.100 163.400 105.100 ;
        RECT 164.100 104.700 165.000 105.100 ;
        RECT 166.200 104.800 168.200 105.100 ;
        RECT 164.100 101.100 164.500 104.700 ;
        RECT 166.200 101.100 166.600 104.800 ;
        RECT 167.800 101.100 168.200 104.800 ;
        RECT 168.600 101.100 169.000 105.100 ;
        RECT 169.400 104.800 170.700 105.100 ;
        RECT 169.400 101.100 169.800 104.800 ;
        RECT 171.000 104.600 171.500 105.100 ;
        RECT 172.600 105.100 173.000 105.200 ;
        RECT 173.600 105.100 173.900 106.800 ;
        RECT 174.200 106.100 174.600 106.600 ;
        RECT 175.800 106.100 176.200 109.900 ;
        RECT 176.600 108.100 177.000 108.600 ;
        RECT 177.400 108.100 177.800 109.900 ;
        RECT 179.500 109.200 180.100 109.900 ;
        RECT 179.500 108.900 180.200 109.200 ;
        RECT 181.800 108.900 182.200 109.900 ;
        RECT 184.000 109.200 184.400 109.900 ;
        RECT 184.000 108.900 185.000 109.200 ;
        RECT 179.800 108.500 180.200 108.900 ;
        RECT 181.900 108.600 182.200 108.900 ;
        RECT 181.900 108.300 183.300 108.600 ;
        RECT 182.900 108.200 183.300 108.300 ;
        RECT 183.800 108.200 184.200 108.600 ;
        RECT 184.600 108.500 185.000 108.900 ;
        RECT 176.600 107.800 177.800 108.100 ;
        RECT 174.200 105.800 176.200 106.100 ;
        RECT 172.600 104.800 173.300 105.100 ;
        RECT 173.600 104.800 174.100 105.100 ;
        RECT 171.000 101.100 171.400 104.600 ;
        RECT 173.000 104.200 173.300 104.800 ;
        RECT 173.000 103.800 173.400 104.200 ;
        RECT 173.700 101.100 174.100 104.800 ;
        RECT 175.800 101.100 176.200 105.800 ;
        RECT 177.400 107.700 177.800 107.800 ;
        RECT 178.900 107.700 179.300 107.800 ;
        RECT 177.400 107.400 179.300 107.700 ;
        RECT 177.400 105.700 177.800 107.400 ;
        RECT 180.900 107.100 181.300 107.200 ;
        RECT 183.800 107.100 184.100 108.200 ;
        RECT 186.200 107.500 186.600 109.900 ;
        RECT 187.000 108.500 187.400 109.500 ;
        RECT 187.000 107.400 187.300 108.500 ;
        RECT 189.100 108.000 189.500 109.500 ;
        RECT 191.800 108.500 192.200 109.500 ;
        RECT 189.100 107.700 189.900 108.000 ;
        RECT 189.500 107.500 189.900 107.700 ;
        RECT 185.400 107.100 186.200 107.200 ;
        RECT 187.000 107.100 189.100 107.400 ;
        RECT 180.700 106.800 186.200 107.100 ;
        RECT 188.600 106.900 189.100 107.100 ;
        RECT 189.600 107.200 189.900 107.500 ;
        RECT 191.800 107.400 192.100 108.500 ;
        RECT 193.900 108.000 194.300 109.500 ;
        RECT 196.600 108.000 197.000 109.900 ;
        RECT 198.200 108.000 198.600 109.900 ;
        RECT 193.900 107.700 194.700 108.000 ;
        RECT 196.600 107.900 198.600 108.000 ;
        RECT 199.000 107.900 199.400 109.900 ;
        RECT 200.100 108.200 200.500 109.900 ;
        RECT 202.500 108.200 202.900 109.900 ;
        RECT 200.100 107.900 201.000 108.200 ;
        RECT 202.500 107.900 203.400 108.200 ;
        RECT 196.700 107.700 198.500 107.900 ;
        RECT 194.300 107.500 194.700 107.700 ;
        RECT 179.800 106.400 180.200 106.500 ;
        RECT 178.300 106.100 180.200 106.400 ;
        RECT 178.300 106.000 178.700 106.100 ;
        RECT 179.100 105.700 179.500 105.800 ;
        RECT 177.400 105.400 179.500 105.700 ;
        RECT 177.400 101.100 177.800 105.400 ;
        RECT 180.700 105.200 181.000 106.800 ;
        RECT 184.300 106.700 184.700 106.800 ;
        RECT 183.800 106.200 184.200 106.300 ;
        RECT 185.100 106.200 185.500 106.300 ;
        RECT 183.000 105.900 185.500 106.200 ;
        RECT 183.000 105.800 183.400 105.900 ;
        RECT 187.000 105.800 187.400 106.600 ;
        RECT 187.800 105.800 188.200 106.600 ;
        RECT 188.600 106.500 189.300 106.900 ;
        RECT 189.600 106.800 190.600 107.200 ;
        RECT 191.800 107.100 193.900 107.400 ;
        RECT 193.400 106.900 193.900 107.100 ;
        RECT 194.400 107.200 194.700 107.500 ;
        RECT 197.000 107.200 197.400 107.400 ;
        RECT 199.000 107.200 199.300 107.900 ;
        RECT 183.800 105.500 186.600 105.600 ;
        RECT 188.600 105.500 188.900 106.500 ;
        RECT 183.700 105.400 186.600 105.500 ;
        RECT 179.800 104.900 181.000 105.200 ;
        RECT 181.700 105.300 186.600 105.400 ;
        RECT 181.700 105.100 184.100 105.300 ;
        RECT 179.800 104.400 180.100 104.900 ;
        RECT 179.400 104.000 180.100 104.400 ;
        RECT 180.900 104.500 181.300 104.600 ;
        RECT 181.700 104.500 182.000 105.100 ;
        RECT 180.900 104.200 182.000 104.500 ;
        RECT 182.300 104.500 185.000 104.800 ;
        RECT 182.300 104.400 182.700 104.500 ;
        RECT 184.600 104.400 185.000 104.500 ;
        RECT 181.500 103.700 181.900 103.800 ;
        RECT 182.900 103.700 183.300 103.800 ;
        RECT 179.800 103.100 180.200 103.500 ;
        RECT 181.500 103.400 183.300 103.700 ;
        RECT 181.900 103.100 182.200 103.400 ;
        RECT 184.600 103.100 185.000 103.500 ;
        RECT 179.500 101.100 180.100 103.100 ;
        RECT 181.800 101.100 182.200 103.100 ;
        RECT 184.000 102.800 185.000 103.100 ;
        RECT 184.000 101.100 184.400 102.800 ;
        RECT 186.200 101.100 186.600 105.300 ;
        RECT 187.000 105.200 188.900 105.500 ;
        RECT 187.000 103.500 187.300 105.200 ;
        RECT 189.600 104.900 189.900 106.800 ;
        RECT 190.200 105.400 190.600 106.200 ;
        RECT 191.800 105.800 192.200 106.600 ;
        RECT 192.600 105.800 193.000 106.600 ;
        RECT 193.400 106.500 194.100 106.900 ;
        RECT 194.400 106.800 195.400 107.200 ;
        RECT 196.600 106.900 197.400 107.200 ;
        RECT 196.600 106.800 197.000 106.900 ;
        RECT 198.100 106.800 199.400 107.200 ;
        RECT 193.400 105.500 193.700 106.500 ;
        RECT 189.100 104.600 189.900 104.900 ;
        RECT 191.800 105.200 193.700 105.500 ;
        RECT 194.400 105.200 194.700 106.800 ;
        RECT 195.000 106.100 195.400 106.200 ;
        RECT 195.800 106.100 196.200 106.200 ;
        RECT 195.000 105.800 196.200 106.100 ;
        RECT 196.600 106.100 197.000 106.200 ;
        RECT 197.400 106.100 197.800 106.600 ;
        RECT 196.600 105.800 197.800 106.100 ;
        RECT 195.000 105.400 195.400 105.800 ;
        RECT 187.000 101.500 187.400 103.500 ;
        RECT 189.100 102.200 189.500 104.600 ;
        RECT 191.800 103.500 192.100 105.200 ;
        RECT 194.200 104.900 194.700 105.200 ;
        RECT 198.100 105.100 198.400 106.800 ;
        RECT 200.600 106.100 201.000 107.900 ;
        RECT 201.400 106.800 201.800 107.600 ;
        RECT 199.000 105.800 201.000 106.100 ;
        RECT 199.000 105.200 199.300 105.800 ;
        RECT 199.000 105.100 199.400 105.200 ;
        RECT 193.900 104.600 194.700 104.900 ;
        RECT 197.900 104.800 198.400 105.100 ;
        RECT 198.700 104.800 199.400 105.100 ;
        RECT 189.100 101.800 189.800 102.200 ;
        RECT 189.100 101.100 189.500 101.800 ;
        RECT 191.800 101.500 192.200 103.500 ;
        RECT 193.900 101.100 194.300 104.600 ;
        RECT 197.900 101.100 198.300 104.800 ;
        RECT 198.700 104.200 199.000 104.800 ;
        RECT 199.800 104.400 200.200 105.200 ;
        RECT 198.600 103.800 199.000 104.200 ;
        RECT 200.600 101.100 201.000 105.800 ;
        RECT 202.200 104.400 202.600 105.200 ;
        RECT 203.000 101.100 203.400 107.900 ;
        RECT 1.400 95.600 1.800 99.900 ;
        RECT 3.000 95.600 3.400 99.900 ;
        RECT 4.600 95.600 5.000 99.900 ;
        RECT 6.200 95.600 6.600 99.900 ;
        RECT 7.800 95.700 8.200 99.900 ;
        RECT 10.000 98.200 10.400 99.900 ;
        RECT 9.400 97.900 10.400 98.200 ;
        RECT 12.200 97.900 12.600 99.900 ;
        RECT 14.300 97.900 14.900 99.900 ;
        RECT 9.400 97.500 9.800 97.900 ;
        RECT 12.200 97.600 12.500 97.900 ;
        RECT 11.100 97.300 12.900 97.600 ;
        RECT 14.200 97.500 14.600 97.900 ;
        RECT 11.100 97.200 11.500 97.300 ;
        RECT 12.500 97.200 12.900 97.300 ;
        RECT 9.400 96.500 9.800 96.600 ;
        RECT 11.700 96.500 12.100 96.600 ;
        RECT 9.400 96.200 12.100 96.500 ;
        RECT 12.400 96.500 13.500 96.800 ;
        RECT 12.400 95.900 12.700 96.500 ;
        RECT 13.100 96.400 13.500 96.500 ;
        RECT 14.300 96.600 15.000 97.000 ;
        RECT 14.300 96.100 14.600 96.600 ;
        RECT 10.300 95.700 12.700 95.900 ;
        RECT 7.800 95.600 12.700 95.700 ;
        RECT 13.400 95.800 14.600 96.100 ;
        RECT 1.400 95.200 2.300 95.600 ;
        RECT 3.000 95.200 4.100 95.600 ;
        RECT 4.600 95.200 5.700 95.600 ;
        RECT 6.200 95.200 7.400 95.600 ;
        RECT 7.800 95.500 10.700 95.600 ;
        RECT 7.800 95.400 10.600 95.500 ;
        RECT 1.900 94.500 2.300 95.200 ;
        RECT 3.700 94.500 4.100 95.200 ;
        RECT 5.300 94.500 5.700 95.200 ;
        RECT 1.900 94.100 3.200 94.500 ;
        RECT 3.700 94.100 4.900 94.500 ;
        RECT 5.300 94.100 6.600 94.500 ;
        RECT 1.900 93.800 2.300 94.100 ;
        RECT 3.700 93.800 4.100 94.100 ;
        RECT 5.300 93.800 5.700 94.100 ;
        RECT 7.000 93.800 7.400 95.200 ;
        RECT 11.000 95.100 11.400 95.200 ;
        RECT 11.800 95.100 12.200 95.200 ;
        RECT 8.900 94.800 12.200 95.100 ;
        RECT 8.900 94.700 9.300 94.800 ;
        RECT 9.700 94.200 10.100 94.300 ;
        RECT 13.400 94.200 13.700 95.800 ;
        RECT 16.600 95.600 17.000 99.900 ;
        RECT 18.700 96.200 19.100 99.900 ;
        RECT 19.400 96.800 19.800 97.200 ;
        RECT 19.500 96.200 19.800 96.800 ;
        RECT 18.700 95.900 19.200 96.200 ;
        RECT 19.500 96.100 20.200 96.200 ;
        RECT 21.400 96.100 21.800 99.900 ;
        RECT 19.500 95.900 21.800 96.100 ;
        RECT 14.900 95.300 17.000 95.600 ;
        RECT 14.900 95.200 15.300 95.300 ;
        RECT 15.700 94.900 16.100 95.000 ;
        RECT 14.200 94.600 16.100 94.900 ;
        RECT 14.200 94.500 14.600 94.600 ;
        RECT 8.200 93.900 13.700 94.200 ;
        RECT 8.200 93.800 9.000 93.900 ;
        RECT 1.400 93.400 2.300 93.800 ;
        RECT 3.000 93.400 4.100 93.800 ;
        RECT 4.600 93.400 5.700 93.800 ;
        RECT 6.200 93.400 7.400 93.800 ;
        RECT 1.400 91.100 1.800 93.400 ;
        RECT 3.000 91.100 3.400 93.400 ;
        RECT 4.600 91.100 5.000 93.400 ;
        RECT 6.200 91.100 6.600 93.400 ;
        RECT 7.800 91.100 8.200 93.500 ;
        RECT 10.300 92.800 10.600 93.900 ;
        RECT 13.100 93.800 13.500 93.900 ;
        RECT 16.600 93.600 17.000 95.300 ;
        RECT 18.900 95.200 19.200 95.900 ;
        RECT 19.800 95.800 21.800 95.900 ;
        RECT 22.200 95.800 22.600 96.600 ;
        RECT 23.000 96.200 23.400 99.900 ;
        RECT 24.600 96.200 25.000 99.900 ;
        RECT 23.000 95.900 25.000 96.200 ;
        RECT 25.400 95.900 25.800 99.900 ;
        RECT 18.200 94.400 18.600 95.200 ;
        RECT 18.900 94.800 19.400 95.200 ;
        RECT 18.900 94.200 19.200 94.800 ;
        RECT 17.400 94.100 17.800 94.200 ;
        RECT 17.400 93.800 18.200 94.100 ;
        RECT 18.900 93.800 20.200 94.200 ;
        RECT 17.800 93.600 18.200 93.800 ;
        RECT 15.100 93.300 17.000 93.600 ;
        RECT 15.100 93.200 15.500 93.300 ;
        RECT 9.400 92.100 9.800 92.500 ;
        RECT 10.200 92.400 10.600 92.800 ;
        RECT 11.100 92.700 11.500 92.800 ;
        RECT 11.100 92.400 12.500 92.700 ;
        RECT 12.200 92.100 12.500 92.400 ;
        RECT 14.200 92.100 14.600 92.500 ;
        RECT 9.400 91.800 10.400 92.100 ;
        RECT 10.000 91.100 10.400 91.800 ;
        RECT 12.200 91.100 12.600 92.100 ;
        RECT 14.200 91.800 14.900 92.100 ;
        RECT 14.300 91.100 14.900 91.800 ;
        RECT 16.600 91.100 17.000 93.300 ;
        RECT 17.500 93.100 19.300 93.300 ;
        RECT 19.800 93.100 20.100 93.800 ;
        RECT 20.600 93.400 21.000 94.200 ;
        RECT 21.400 93.100 21.800 95.800 ;
        RECT 23.400 95.200 23.800 95.400 ;
        RECT 25.400 95.200 25.700 95.900 ;
        RECT 22.200 95.100 22.600 95.200 ;
        RECT 23.000 95.100 23.800 95.200 ;
        RECT 22.200 94.900 23.800 95.100 ;
        RECT 24.600 94.900 25.800 95.200 ;
        RECT 22.200 94.800 23.400 94.900 ;
        RECT 23.800 93.800 24.200 94.600 ;
        RECT 24.600 93.100 24.900 94.900 ;
        RECT 25.400 94.800 25.800 94.900 ;
        RECT 17.400 93.000 19.400 93.100 ;
        RECT 17.400 91.100 17.800 93.000 ;
        RECT 19.000 91.100 19.400 93.000 ;
        RECT 19.800 91.100 20.200 93.100 ;
        RECT 21.400 92.800 22.300 93.100 ;
        RECT 21.900 91.100 22.300 92.800 ;
        RECT 24.600 91.100 25.000 93.100 ;
        RECT 25.400 92.800 25.800 93.200 ;
        RECT 25.300 92.400 25.700 92.800 ;
        RECT 26.200 92.400 26.600 93.200 ;
        RECT 27.000 91.100 27.400 99.900 ;
        RECT 27.800 96.200 28.200 99.900 ;
        RECT 29.400 96.200 29.800 99.900 ;
        RECT 27.800 95.900 29.800 96.200 ;
        RECT 30.200 95.900 30.600 99.900 ;
        RECT 31.000 96.200 31.400 99.900 ;
        RECT 32.600 96.200 33.000 99.900 ;
        RECT 31.000 95.900 33.000 96.200 ;
        RECT 33.400 95.900 33.800 99.900 ;
        RECT 35.500 96.200 35.900 99.900 ;
        RECT 36.200 96.800 36.600 97.200 ;
        RECT 36.300 96.200 36.600 96.800 ;
        RECT 38.700 96.200 39.100 99.900 ;
        RECT 39.400 96.800 39.800 97.200 ;
        RECT 39.500 96.200 39.800 96.800 ;
        RECT 35.500 95.900 36.000 96.200 ;
        RECT 36.300 95.900 37.000 96.200 ;
        RECT 38.700 95.900 39.200 96.200 ;
        RECT 39.500 95.900 40.200 96.200 ;
        RECT 40.600 95.900 41.000 99.900 ;
        RECT 41.400 96.200 41.800 99.900 ;
        RECT 43.000 96.200 43.400 99.900 ;
        RECT 44.200 96.800 44.600 97.200 ;
        RECT 44.200 96.200 44.500 96.800 ;
        RECT 44.900 96.200 45.300 99.900 ;
        RECT 41.400 95.900 43.400 96.200 ;
        RECT 43.800 95.900 44.500 96.200 ;
        RECT 44.800 95.900 45.300 96.200 ;
        RECT 48.300 95.900 49.300 99.900 ;
        RECT 53.400 96.400 53.800 99.900 ;
        RECT 53.300 95.900 53.800 96.400 ;
        RECT 55.000 96.200 55.400 99.900 ;
        RECT 56.200 96.800 56.600 97.200 ;
        RECT 56.200 96.200 56.500 96.800 ;
        RECT 56.900 96.200 57.300 99.900 ;
        RECT 59.000 96.200 59.400 99.900 ;
        RECT 60.600 96.200 61.000 99.900 ;
        RECT 54.100 95.900 55.400 96.200 ;
        RECT 55.800 95.900 56.500 96.200 ;
        RECT 28.200 95.200 28.600 95.400 ;
        RECT 30.200 95.200 30.500 95.900 ;
        RECT 31.400 95.200 31.800 95.400 ;
        RECT 33.400 95.200 33.700 95.900 ;
        RECT 27.800 94.900 28.600 95.200 ;
        RECT 29.400 94.900 30.600 95.200 ;
        RECT 27.800 94.800 28.200 94.900 ;
        RECT 27.800 94.100 28.200 94.200 ;
        RECT 28.600 94.100 29.000 94.600 ;
        RECT 27.800 93.800 29.000 94.100 ;
        RECT 29.400 93.100 29.700 94.900 ;
        RECT 30.200 94.800 30.600 94.900 ;
        RECT 31.000 94.900 31.800 95.200 ;
        RECT 32.600 95.100 33.800 95.200 ;
        RECT 34.200 95.100 34.600 95.200 ;
        RECT 32.600 94.900 34.600 95.100 ;
        RECT 31.000 94.800 31.400 94.900 ;
        RECT 31.800 93.800 32.200 94.600 ;
        RECT 29.400 91.100 29.800 93.100 ;
        RECT 30.200 92.800 30.600 93.200 ;
        RECT 32.600 93.100 32.900 94.900 ;
        RECT 33.400 94.800 34.600 94.900 ;
        RECT 35.000 94.400 35.400 95.200 ;
        RECT 35.700 94.200 36.000 95.900 ;
        RECT 36.600 95.800 37.000 95.900 ;
        RECT 37.400 95.100 37.800 95.200 ;
        RECT 38.200 95.100 38.600 95.200 ;
        RECT 37.400 94.800 38.600 95.100 ;
        RECT 38.200 94.400 38.600 94.800 ;
        RECT 38.900 94.200 39.200 95.900 ;
        RECT 39.800 95.800 40.200 95.900 ;
        RECT 40.700 95.200 41.000 95.900 ;
        RECT 43.800 95.800 44.200 95.900 ;
        RECT 42.600 95.200 43.000 95.400 ;
        RECT 40.600 94.900 41.800 95.200 ;
        RECT 42.600 94.900 43.400 95.200 ;
        RECT 40.600 94.800 41.000 94.900 ;
        RECT 41.400 94.800 41.800 94.900 ;
        RECT 43.000 94.800 43.400 94.900 ;
        RECT 34.200 94.100 34.600 94.200 ;
        RECT 34.200 93.800 35.000 94.100 ;
        RECT 35.700 93.800 37.000 94.200 ;
        RECT 37.400 94.100 37.800 94.200 ;
        RECT 37.400 93.800 38.200 94.100 ;
        RECT 38.900 93.800 40.200 94.200 ;
        RECT 34.600 93.600 35.000 93.800 ;
        RECT 30.100 92.400 30.500 92.800 ;
        RECT 32.600 91.100 33.000 93.100 ;
        RECT 33.400 92.800 33.800 93.200 ;
        RECT 34.300 93.100 36.100 93.300 ;
        RECT 36.600 93.100 36.900 93.800 ;
        RECT 37.800 93.600 38.200 93.800 ;
        RECT 37.500 93.100 39.300 93.300 ;
        RECT 39.800 93.100 40.100 93.800 ;
        RECT 40.600 93.100 41.000 93.200 ;
        RECT 41.500 93.100 41.800 94.800 ;
        RECT 42.200 93.800 42.600 94.600 ;
        RECT 44.800 94.200 45.100 95.900 ;
        RECT 45.400 94.400 45.800 95.200 ;
        RECT 47.800 94.400 48.200 95.200 ;
        RECT 48.600 94.200 48.900 95.900 ;
        RECT 49.400 94.400 49.800 95.200 ;
        RECT 43.800 93.800 45.100 94.200 ;
        RECT 46.200 94.100 46.600 94.200 ;
        RECT 45.800 93.800 46.600 94.100 ;
        RECT 47.000 94.100 47.400 94.200 ;
        RECT 48.600 94.100 49.000 94.200 ;
        RECT 50.200 94.100 50.600 94.600 ;
        RECT 53.300 94.200 53.600 95.900 ;
        RECT 54.100 94.900 54.400 95.900 ;
        RECT 55.800 95.800 56.200 95.900 ;
        RECT 56.800 95.800 57.800 96.200 ;
        RECT 59.000 95.900 61.000 96.200 ;
        RECT 61.400 95.900 61.800 99.900 ;
        RECT 62.200 95.900 62.600 99.900 ;
        RECT 63.000 96.200 63.400 99.900 ;
        RECT 64.600 96.200 65.000 99.900 ;
        RECT 63.000 95.900 65.000 96.200 ;
        RECT 65.400 96.200 65.800 99.900 ;
        RECT 67.000 96.400 67.400 99.900 ;
        RECT 65.400 95.900 66.700 96.200 ;
        RECT 67.000 95.900 67.500 96.400 ;
        RECT 53.900 94.500 54.400 94.900 ;
        RECT 51.000 94.100 51.400 94.200 ;
        RECT 47.000 93.800 47.800 94.100 ;
        RECT 48.600 93.800 49.800 94.100 ;
        RECT 50.200 93.800 51.400 94.100 ;
        RECT 53.300 93.800 53.800 94.200 ;
        RECT 43.900 93.100 44.200 93.800 ;
        RECT 45.800 93.600 46.200 93.800 ;
        RECT 47.400 93.600 47.800 93.800 ;
        RECT 44.700 93.100 46.500 93.300 ;
        RECT 47.100 93.100 48.900 93.300 ;
        RECT 49.500 93.100 49.800 93.800 ;
        RECT 53.300 93.200 53.600 93.800 ;
        RECT 54.100 93.700 54.400 94.500 ;
        RECT 54.900 95.100 55.400 95.200 ;
        RECT 55.800 95.100 56.200 95.200 ;
        RECT 54.900 94.800 56.200 95.100 ;
        RECT 54.900 94.400 55.300 94.800 ;
        RECT 56.800 94.200 57.100 95.800 ;
        RECT 59.400 95.200 59.800 95.400 ;
        RECT 61.400 95.200 61.700 95.900 ;
        RECT 62.300 95.200 62.600 95.900 ;
        RECT 64.200 95.200 64.600 95.400 ;
        RECT 57.400 94.400 57.800 95.200 ;
        RECT 58.200 95.100 58.600 95.200 ;
        RECT 59.000 95.100 59.800 95.200 ;
        RECT 58.200 94.900 59.800 95.100 ;
        RECT 60.600 94.900 61.800 95.200 ;
        RECT 58.200 94.800 59.400 94.900 ;
        RECT 55.800 93.800 57.100 94.200 ;
        RECT 58.200 94.100 58.600 94.200 ;
        RECT 57.800 93.800 58.600 94.100 ;
        RECT 59.800 93.800 60.200 94.600 ;
        RECT 60.600 94.100 60.900 94.900 ;
        RECT 61.400 94.800 61.800 94.900 ;
        RECT 62.200 94.900 63.400 95.200 ;
        RECT 64.200 94.900 65.000 95.200 ;
        RECT 62.200 94.800 62.600 94.900 ;
        RECT 60.600 93.800 62.500 94.100 ;
        RECT 54.100 93.400 55.400 93.700 ;
        RECT 34.200 93.000 36.200 93.100 ;
        RECT 33.300 92.400 33.700 92.800 ;
        RECT 34.200 91.100 34.600 93.000 ;
        RECT 35.800 91.100 36.200 93.000 ;
        RECT 36.600 91.100 37.000 93.100 ;
        RECT 37.400 93.000 39.400 93.100 ;
        RECT 37.400 91.100 37.800 93.000 ;
        RECT 39.000 91.100 39.400 93.000 ;
        RECT 39.800 92.800 41.000 93.100 ;
        RECT 39.800 91.100 40.200 92.800 ;
        RECT 40.700 92.400 41.100 92.800 ;
        RECT 41.400 91.100 41.800 93.100 ;
        RECT 43.800 91.100 44.200 93.100 ;
        RECT 44.600 93.000 46.600 93.100 ;
        RECT 44.600 91.100 45.000 93.000 ;
        RECT 46.200 91.100 46.600 93.000 ;
        RECT 47.000 93.000 49.000 93.100 ;
        RECT 47.000 91.100 47.400 93.000 ;
        RECT 48.600 91.400 49.000 93.000 ;
        RECT 49.400 91.700 49.800 93.100 ;
        RECT 50.200 91.400 50.600 93.100 ;
        RECT 53.300 92.800 53.800 93.200 ;
        RECT 48.600 91.100 50.600 91.400 ;
        RECT 53.400 91.100 53.800 92.800 ;
        RECT 55.000 91.100 55.400 93.400 ;
        RECT 55.900 93.100 56.200 93.800 ;
        RECT 57.800 93.600 58.200 93.800 ;
        RECT 56.700 93.100 58.500 93.300 ;
        RECT 60.600 93.100 60.900 93.800 ;
        RECT 62.200 93.200 62.500 93.800 ;
        RECT 55.800 91.100 56.200 93.100 ;
        RECT 56.600 93.000 58.600 93.100 ;
        RECT 56.600 91.100 57.000 93.000 ;
        RECT 58.200 91.100 58.600 93.000 ;
        RECT 60.600 91.100 61.000 93.100 ;
        RECT 61.400 92.800 61.800 93.200 ;
        RECT 62.200 92.800 62.600 93.200 ;
        RECT 63.100 93.100 63.400 94.900 ;
        RECT 64.600 94.800 65.000 94.900 ;
        RECT 65.400 94.800 65.900 95.200 ;
        RECT 63.800 93.800 64.200 94.600 ;
        RECT 65.500 94.400 65.900 94.800 ;
        RECT 66.400 94.900 66.700 95.900 ;
        RECT 66.400 94.500 66.900 94.900 ;
        RECT 66.400 93.700 66.700 94.500 ;
        RECT 67.200 94.200 67.500 95.900 ;
        RECT 67.000 93.800 67.500 94.200 ;
        RECT 61.300 92.400 61.700 92.800 ;
        RECT 62.300 92.400 62.700 92.800 ;
        RECT 63.000 91.100 63.400 93.100 ;
        RECT 65.400 93.400 66.700 93.700 ;
        RECT 65.400 91.100 65.800 93.400 ;
        RECT 67.200 93.100 67.500 93.800 ;
        RECT 67.000 92.800 67.500 93.100 ;
        RECT 69.400 95.600 69.800 99.900 ;
        RECT 71.000 95.600 71.400 99.900 ;
        RECT 73.900 95.900 74.900 99.900 ;
        RECT 77.000 96.800 77.400 97.200 ;
        RECT 77.000 96.200 77.300 96.800 ;
        RECT 77.700 96.200 78.100 99.900 ;
        RECT 80.900 98.200 81.300 99.900 ;
        RECT 80.900 97.800 81.800 98.200 ;
        RECT 80.200 96.800 80.600 97.200 ;
        RECT 80.200 96.200 80.500 96.800 ;
        RECT 80.900 96.200 81.300 97.800 ;
        RECT 83.400 96.800 83.800 97.200 ;
        RECT 83.400 96.200 83.700 96.800 ;
        RECT 84.100 96.200 84.500 99.900 ;
        RECT 76.600 95.900 77.300 96.200 ;
        RECT 77.600 95.900 78.100 96.200 ;
        RECT 79.800 95.900 80.500 96.200 ;
        RECT 80.800 95.900 81.300 96.200 ;
        RECT 83.000 95.900 83.700 96.200 ;
        RECT 84.000 95.900 84.500 96.200 ;
        RECT 87.500 95.900 88.500 99.900 ;
        RECT 90.200 95.900 90.600 99.900 ;
        RECT 91.000 96.200 91.400 99.900 ;
        RECT 92.600 96.200 93.000 99.900 ;
        RECT 93.800 96.800 94.200 97.200 ;
        RECT 93.800 96.200 94.100 96.800 ;
        RECT 94.500 96.200 94.900 99.900 ;
        RECT 97.400 96.400 97.800 99.900 ;
        RECT 91.000 95.900 93.000 96.200 ;
        RECT 93.400 95.900 94.100 96.200 ;
        RECT 94.400 95.900 94.900 96.200 ;
        RECT 97.300 95.900 97.800 96.400 ;
        RECT 99.000 96.200 99.400 99.900 ;
        RECT 100.600 96.400 101.000 99.900 ;
        RECT 98.100 95.900 99.400 96.200 ;
        RECT 100.500 95.900 101.000 96.400 ;
        RECT 102.200 96.200 102.600 99.900 ;
        RECT 101.300 95.900 102.600 96.200 ;
        RECT 69.400 95.200 71.400 95.600 ;
        RECT 74.300 95.200 74.600 95.900 ;
        RECT 76.600 95.800 77.000 95.900 ;
        RECT 69.400 93.800 69.800 95.200 ;
        RECT 69.400 93.400 71.400 93.800 ;
        RECT 71.800 93.400 72.200 94.200 ;
        RECT 72.600 93.800 73.000 94.600 ;
        RECT 73.400 94.400 73.800 95.200 ;
        RECT 74.200 94.800 74.600 95.200 ;
        RECT 74.300 94.200 74.600 94.800 ;
        RECT 75.000 94.400 75.400 95.200 ;
        RECT 75.800 95.100 76.200 95.200 ;
        RECT 77.600 95.100 77.900 95.900 ;
        RECT 79.800 95.800 80.200 95.900 ;
        RECT 75.800 94.800 77.900 95.100 ;
        RECT 77.600 94.200 77.900 94.800 ;
        RECT 78.200 94.400 78.600 95.200 ;
        RECT 80.800 94.200 81.100 95.900 ;
        RECT 83.000 95.800 83.400 95.900 ;
        RECT 81.400 95.100 81.800 95.200 ;
        RECT 83.000 95.100 83.400 95.200 ;
        RECT 81.400 94.800 83.400 95.100 ;
        RECT 81.400 94.400 81.800 94.800 ;
        RECT 84.000 94.200 84.300 95.900 ;
        RECT 84.600 94.400 85.000 95.200 ;
        RECT 87.000 94.400 87.400 95.200 ;
        RECT 87.800 94.200 88.100 95.900 ;
        RECT 90.300 95.200 90.600 95.900 ;
        RECT 93.400 95.800 93.800 95.900 ;
        RECT 92.200 95.200 92.600 95.400 ;
        RECT 88.600 94.400 89.000 95.200 ;
        RECT 90.200 94.900 91.400 95.200 ;
        RECT 92.200 94.900 93.000 95.200 ;
        RECT 90.200 94.800 90.600 94.900 ;
        RECT 74.200 94.100 74.600 94.200 ;
        RECT 75.800 94.100 76.200 94.200 ;
        RECT 73.400 93.800 74.600 94.100 ;
        RECT 75.400 93.800 76.200 94.100 ;
        RECT 76.600 93.800 77.900 94.200 ;
        RECT 79.000 94.100 79.400 94.200 ;
        RECT 78.600 93.800 79.400 94.100 ;
        RECT 79.800 93.800 81.100 94.200 ;
        RECT 82.200 94.100 82.600 94.200 ;
        RECT 81.800 93.800 82.600 94.100 ;
        RECT 83.000 93.800 84.300 94.200 ;
        RECT 85.400 94.100 85.800 94.200 ;
        RECT 85.000 93.800 85.800 94.100 ;
        RECT 86.200 94.100 86.600 94.200 ;
        RECT 87.800 94.100 88.200 94.200 ;
        RECT 89.400 94.100 89.800 94.600 ;
        RECT 90.200 94.100 90.600 94.200 ;
        RECT 86.200 93.800 87.000 94.100 ;
        RECT 87.800 93.800 89.000 94.100 ;
        RECT 89.400 93.800 90.600 94.100 ;
        RECT 67.000 91.100 67.400 92.800 ;
        RECT 69.400 91.100 69.800 93.400 ;
        RECT 71.000 91.100 71.400 93.400 ;
        RECT 73.400 93.100 73.700 93.800 ;
        RECT 75.400 93.600 75.800 93.800 ;
        RECT 74.300 93.100 76.100 93.300 ;
        RECT 76.700 93.100 77.000 93.800 ;
        RECT 78.600 93.600 79.000 93.800 ;
        RECT 77.500 93.100 79.300 93.300 ;
        RECT 79.900 93.100 80.200 93.800 ;
        RECT 81.800 93.600 82.200 93.800 ;
        RECT 80.700 93.100 82.500 93.300 ;
        RECT 83.100 93.200 83.400 93.800 ;
        RECT 85.000 93.600 85.400 93.800 ;
        RECT 86.600 93.600 87.000 93.800 ;
        RECT 72.600 91.400 73.000 93.100 ;
        RECT 73.400 91.700 73.800 93.100 ;
        RECT 74.200 93.000 76.200 93.100 ;
        RECT 74.200 91.400 74.600 93.000 ;
        RECT 72.600 91.100 74.600 91.400 ;
        RECT 75.800 91.100 76.200 93.000 ;
        RECT 76.600 91.100 77.000 93.100 ;
        RECT 77.400 93.000 79.400 93.100 ;
        RECT 77.400 91.100 77.800 93.000 ;
        RECT 79.000 91.100 79.400 93.000 ;
        RECT 79.800 91.100 80.200 93.100 ;
        RECT 80.600 93.000 82.600 93.100 ;
        RECT 80.600 91.100 81.000 93.000 ;
        RECT 82.200 91.100 82.600 93.000 ;
        RECT 83.000 91.100 83.400 93.200 ;
        RECT 83.900 93.100 85.700 93.300 ;
        RECT 86.300 93.100 88.100 93.300 ;
        RECT 88.700 93.100 89.000 93.800 ;
        RECT 83.800 93.000 85.800 93.100 ;
        RECT 83.800 91.100 84.200 93.000 ;
        RECT 85.400 91.100 85.800 93.000 ;
        RECT 86.200 93.000 88.200 93.100 ;
        RECT 86.200 91.100 86.600 93.000 ;
        RECT 87.800 91.400 88.200 93.000 ;
        RECT 88.600 91.700 89.000 93.100 ;
        RECT 89.400 91.400 89.800 93.100 ;
        RECT 90.200 92.800 90.600 93.200 ;
        RECT 91.100 93.100 91.400 94.900 ;
        RECT 92.600 94.800 93.000 94.900 ;
        RECT 91.800 93.800 92.200 94.600 ;
        RECT 94.400 94.200 94.700 95.900 ;
        RECT 95.000 95.100 95.400 95.200 ;
        RECT 95.800 95.100 96.200 95.200 ;
        RECT 95.000 94.800 96.200 95.100 ;
        RECT 95.000 94.400 95.400 94.800 ;
        RECT 97.300 94.200 97.600 95.900 ;
        RECT 98.100 94.900 98.400 95.900 ;
        RECT 97.900 94.500 98.400 94.900 ;
        RECT 93.400 93.800 94.700 94.200 ;
        RECT 95.800 94.100 96.200 94.200 ;
        RECT 96.600 94.100 97.000 94.200 ;
        RECT 95.400 93.800 97.000 94.100 ;
        RECT 97.300 93.800 97.800 94.200 ;
        RECT 93.500 93.100 93.800 93.800 ;
        RECT 95.400 93.600 95.800 93.800 ;
        RECT 94.300 93.100 96.100 93.300 ;
        RECT 97.300 93.100 97.600 93.800 ;
        RECT 98.100 93.700 98.400 94.500 ;
        RECT 98.900 94.800 99.400 95.200 ;
        RECT 98.900 94.400 99.300 94.800 ;
        RECT 100.500 94.200 100.800 95.900 ;
        RECT 101.300 94.900 101.600 95.900 ;
        RECT 104.600 95.700 105.000 99.900 ;
        RECT 106.800 98.200 107.200 99.900 ;
        RECT 106.200 97.900 107.200 98.200 ;
        RECT 109.000 97.900 109.400 99.900 ;
        RECT 111.100 97.900 111.700 99.900 ;
        RECT 106.200 97.500 106.600 97.900 ;
        RECT 109.000 97.600 109.300 97.900 ;
        RECT 107.900 97.300 109.700 97.600 ;
        RECT 111.000 97.500 111.400 97.900 ;
        RECT 107.900 97.200 108.300 97.300 ;
        RECT 109.300 97.200 109.700 97.300 ;
        RECT 106.200 96.500 106.600 96.600 ;
        RECT 108.500 96.500 108.900 96.600 ;
        RECT 106.200 96.200 108.900 96.500 ;
        RECT 109.200 96.500 110.300 96.800 ;
        RECT 109.200 95.900 109.500 96.500 ;
        RECT 109.900 96.400 110.300 96.500 ;
        RECT 111.100 96.600 111.800 97.000 ;
        RECT 111.100 96.100 111.400 96.600 ;
        RECT 107.100 95.700 109.500 95.900 ;
        RECT 104.600 95.600 109.500 95.700 ;
        RECT 110.200 95.800 111.400 96.100 ;
        RECT 104.600 95.500 107.500 95.600 ;
        RECT 104.600 95.400 107.400 95.500 ;
        RECT 110.200 95.200 110.500 95.800 ;
        RECT 113.400 95.600 113.800 99.900 ;
        RECT 115.500 96.200 115.900 99.900 ;
        RECT 116.200 96.800 116.600 97.200 ;
        RECT 116.300 96.200 116.600 96.800 ;
        RECT 115.500 95.900 116.000 96.200 ;
        RECT 116.300 95.900 117.000 96.200 ;
        RECT 111.700 95.300 113.800 95.600 ;
        RECT 111.700 95.200 112.100 95.300 ;
        RECT 101.100 94.500 101.600 94.900 ;
        RECT 99.800 94.100 100.200 94.200 ;
        RECT 100.500 94.100 101.000 94.200 ;
        RECT 99.800 93.800 101.000 94.100 ;
        RECT 98.100 93.400 99.400 93.700 ;
        RECT 90.300 92.400 90.700 92.800 ;
        RECT 87.800 91.100 89.800 91.400 ;
        RECT 91.000 91.100 91.400 93.100 ;
        RECT 93.400 91.100 93.800 93.100 ;
        RECT 94.200 93.000 96.200 93.100 ;
        RECT 94.200 91.100 94.600 93.000 ;
        RECT 95.800 91.100 96.200 93.000 ;
        RECT 97.300 92.800 97.800 93.100 ;
        RECT 97.400 91.100 97.800 92.800 ;
        RECT 99.000 91.100 99.400 93.400 ;
        RECT 100.500 93.100 100.800 93.800 ;
        RECT 101.300 93.700 101.600 94.500 ;
        RECT 102.100 94.800 102.600 95.200 ;
        RECT 107.800 95.100 108.200 95.200 ;
        RECT 105.700 94.800 108.200 95.100 ;
        RECT 110.200 94.800 110.600 95.200 ;
        RECT 112.500 94.900 112.900 95.000 ;
        RECT 102.100 94.400 102.500 94.800 ;
        RECT 105.700 94.700 106.100 94.800 ;
        RECT 106.500 94.200 106.900 94.300 ;
        RECT 110.200 94.200 110.500 94.800 ;
        RECT 111.000 94.600 112.900 94.900 ;
        RECT 111.000 94.500 111.400 94.600 ;
        RECT 105.000 93.900 110.500 94.200 ;
        RECT 105.000 93.800 105.800 93.900 ;
        RECT 101.300 93.400 102.600 93.700 ;
        RECT 100.500 92.800 101.000 93.100 ;
        RECT 100.600 91.100 101.000 92.800 ;
        RECT 102.200 91.100 102.600 93.400 ;
        RECT 104.600 91.100 105.000 93.500 ;
        RECT 107.100 92.800 107.400 93.900 ;
        RECT 109.900 93.800 110.300 93.900 ;
        RECT 113.400 93.600 113.800 95.300 ;
        RECT 115.000 94.400 115.400 95.200 ;
        RECT 115.700 94.200 116.000 95.900 ;
        RECT 116.600 95.800 117.000 95.900 ;
        RECT 118.200 95.100 118.600 99.900 ;
        RECT 120.200 96.800 120.600 97.200 ;
        RECT 119.000 95.800 119.400 96.600 ;
        RECT 120.200 96.200 120.500 96.800 ;
        RECT 120.900 96.200 121.300 99.900 ;
        RECT 123.800 96.400 124.200 99.900 ;
        RECT 119.800 95.900 120.500 96.200 ;
        RECT 120.800 95.900 121.300 96.200 ;
        RECT 123.700 95.900 124.200 96.400 ;
        RECT 125.400 96.200 125.800 99.900 ;
        RECT 124.500 95.900 125.800 96.200 ;
        RECT 126.200 96.200 126.600 99.900 ;
        RECT 127.800 96.400 128.200 99.900 ;
        RECT 126.200 95.900 127.500 96.200 ;
        RECT 127.800 95.900 128.300 96.400 ;
        RECT 119.800 95.800 120.200 95.900 ;
        RECT 119.800 95.100 120.100 95.800 ;
        RECT 118.200 94.800 120.100 95.100 ;
        RECT 114.200 94.100 114.600 94.200 ;
        RECT 114.200 93.800 115.000 94.100 ;
        RECT 115.700 93.800 117.000 94.200 ;
        RECT 114.600 93.600 115.000 93.800 ;
        RECT 111.900 93.300 113.800 93.600 ;
        RECT 111.900 93.200 112.300 93.300 ;
        RECT 106.200 92.100 106.600 92.500 ;
        RECT 107.000 92.400 107.400 92.800 ;
        RECT 107.900 92.700 108.300 92.800 ;
        RECT 107.900 92.400 109.300 92.700 ;
        RECT 109.000 92.100 109.300 92.400 ;
        RECT 111.000 92.100 111.400 92.500 ;
        RECT 106.200 91.800 107.200 92.100 ;
        RECT 106.800 91.100 107.200 91.800 ;
        RECT 109.000 91.100 109.400 92.100 ;
        RECT 111.000 91.800 111.700 92.100 ;
        RECT 111.100 91.100 111.700 91.800 ;
        RECT 113.400 91.100 113.800 93.300 ;
        RECT 114.300 93.100 116.100 93.300 ;
        RECT 116.600 93.100 116.900 93.800 ;
        RECT 117.400 93.400 117.800 94.200 ;
        RECT 118.200 93.100 118.600 94.800 ;
        RECT 120.800 94.200 121.100 95.900 ;
        RECT 121.400 95.100 121.800 95.200 ;
        RECT 122.200 95.100 122.600 95.200 ;
        RECT 121.400 94.800 122.600 95.100 ;
        RECT 121.400 94.400 121.800 94.800 ;
        RECT 123.700 94.200 124.000 95.900 ;
        RECT 124.500 94.900 124.800 95.900 ;
        RECT 124.300 94.500 124.800 94.900 ;
        RECT 119.000 94.100 119.400 94.200 ;
        RECT 119.800 94.100 121.100 94.200 ;
        RECT 122.200 94.100 122.600 94.200 ;
        RECT 119.000 93.800 121.100 94.100 ;
        RECT 121.800 93.800 122.600 94.100 ;
        RECT 123.700 93.800 124.200 94.200 ;
        RECT 119.900 93.100 120.200 93.800 ;
        RECT 121.800 93.600 122.200 93.800 ;
        RECT 120.700 93.100 122.500 93.300 ;
        RECT 123.700 93.100 124.000 93.800 ;
        RECT 124.500 93.700 124.800 94.500 ;
        RECT 125.300 94.800 125.800 95.200 ;
        RECT 126.200 94.800 126.700 95.200 ;
        RECT 125.300 94.400 125.700 94.800 ;
        RECT 126.300 94.400 126.700 94.800 ;
        RECT 127.200 94.900 127.500 95.900 ;
        RECT 127.200 94.500 127.700 94.900 ;
        RECT 127.200 93.700 127.500 94.500 ;
        RECT 128.000 94.200 128.300 95.900 ;
        RECT 129.400 95.700 129.800 99.900 ;
        RECT 131.600 98.200 132.000 99.900 ;
        RECT 131.000 97.900 132.000 98.200 ;
        RECT 133.800 97.900 134.200 99.900 ;
        RECT 135.900 97.900 136.500 99.900 ;
        RECT 131.000 97.500 131.400 97.900 ;
        RECT 133.800 97.600 134.100 97.900 ;
        RECT 132.700 97.300 134.500 97.600 ;
        RECT 135.800 97.500 136.200 97.900 ;
        RECT 132.700 97.200 133.100 97.300 ;
        RECT 134.100 97.200 134.500 97.300 ;
        RECT 131.000 96.500 131.400 96.600 ;
        RECT 133.300 96.500 133.700 96.600 ;
        RECT 131.000 96.200 133.700 96.500 ;
        RECT 134.000 96.500 135.100 96.800 ;
        RECT 134.000 95.900 134.300 96.500 ;
        RECT 134.700 96.400 135.100 96.500 ;
        RECT 135.900 96.600 136.600 97.000 ;
        RECT 135.900 96.100 136.200 96.600 ;
        RECT 131.900 95.700 134.300 95.900 ;
        RECT 129.400 95.600 134.300 95.700 ;
        RECT 135.000 95.800 136.200 96.100 ;
        RECT 129.400 95.500 132.300 95.600 ;
        RECT 129.400 95.400 132.200 95.500 ;
        RECT 132.600 95.100 133.000 95.200 ;
        RECT 130.500 94.800 133.000 95.100 ;
        RECT 130.500 94.700 130.900 94.800 ;
        RECT 131.300 94.200 131.700 94.300 ;
        RECT 135.000 94.200 135.300 95.800 ;
        RECT 138.200 95.600 138.600 99.900 ;
        RECT 139.000 96.200 139.400 99.900 ;
        RECT 140.600 96.200 141.000 99.900 ;
        RECT 139.000 95.900 141.000 96.200 ;
        RECT 141.400 95.900 141.800 99.900 ;
        RECT 142.500 96.300 142.900 99.900 ;
        RECT 142.500 95.900 143.400 96.300 ;
        RECT 145.900 96.200 146.300 99.900 ;
        RECT 146.600 96.800 147.000 97.200 ;
        RECT 146.700 96.200 147.000 96.800 ;
        RECT 147.800 96.200 148.200 99.900 ;
        RECT 149.400 96.200 149.800 99.900 ;
        RECT 145.900 95.900 146.400 96.200 ;
        RECT 146.700 95.900 147.400 96.200 ;
        RECT 147.800 95.900 149.800 96.200 ;
        RECT 150.200 95.900 150.600 99.900 ;
        RECT 151.000 96.200 151.400 99.900 ;
        RECT 152.600 96.400 153.000 99.900 ;
        RECT 151.000 95.900 152.300 96.200 ;
        RECT 152.600 95.900 153.100 96.400 ;
        RECT 156.100 96.200 156.500 99.900 ;
        RECT 136.500 95.300 138.600 95.600 ;
        RECT 136.500 95.200 136.900 95.300 ;
        RECT 137.300 94.900 137.700 95.000 ;
        RECT 135.800 94.600 137.700 94.900 ;
        RECT 135.800 94.500 136.200 94.600 ;
        RECT 127.800 93.800 128.300 94.200 ;
        RECT 129.800 93.900 135.300 94.200 ;
        RECT 129.800 93.800 130.600 93.900 ;
        RECT 124.500 93.400 125.800 93.700 ;
        RECT 114.200 93.000 116.200 93.100 ;
        RECT 114.200 91.100 114.600 93.000 ;
        RECT 115.800 91.100 116.200 93.000 ;
        RECT 116.600 91.100 117.000 93.100 ;
        RECT 118.200 92.800 119.100 93.100 ;
        RECT 118.700 91.100 119.100 92.800 ;
        RECT 119.800 91.100 120.200 93.100 ;
        RECT 120.600 93.000 122.600 93.100 ;
        RECT 120.600 91.100 121.000 93.000 ;
        RECT 122.200 91.100 122.600 93.000 ;
        RECT 123.700 92.800 124.200 93.100 ;
        RECT 123.800 91.100 124.200 92.800 ;
        RECT 125.400 91.100 125.800 93.400 ;
        RECT 126.200 93.400 127.500 93.700 ;
        RECT 126.200 91.100 126.600 93.400 ;
        RECT 128.000 93.100 128.300 93.800 ;
        RECT 127.800 92.800 128.300 93.100 ;
        RECT 127.800 91.100 128.200 92.800 ;
        RECT 129.400 91.100 129.800 93.500 ;
        RECT 131.900 92.800 132.200 93.900 ;
        RECT 134.700 93.800 135.100 93.900 ;
        RECT 138.200 93.600 138.600 95.300 ;
        RECT 139.400 95.200 139.800 95.400 ;
        RECT 141.400 95.200 141.700 95.900 ;
        RECT 139.000 94.900 139.800 95.200 ;
        RECT 140.600 94.900 141.800 95.200 ;
        RECT 139.000 94.800 139.400 94.900 ;
        RECT 139.800 93.800 140.200 94.600 ;
        RECT 136.700 93.300 138.600 93.600 ;
        RECT 136.700 93.200 137.100 93.300 ;
        RECT 131.000 92.100 131.400 92.500 ;
        RECT 131.800 92.400 132.200 92.800 ;
        RECT 132.700 92.700 133.100 92.800 ;
        RECT 132.700 92.400 134.100 92.700 ;
        RECT 133.800 92.100 134.100 92.400 ;
        RECT 135.800 92.100 136.200 92.500 ;
        RECT 131.000 91.800 132.000 92.100 ;
        RECT 131.600 91.100 132.000 91.800 ;
        RECT 133.800 91.100 134.200 92.100 ;
        RECT 135.800 91.800 136.500 92.100 ;
        RECT 135.900 91.100 136.500 91.800 ;
        RECT 138.200 91.100 138.600 93.300 ;
        RECT 140.600 93.200 140.900 94.900 ;
        RECT 141.400 94.800 141.800 94.900 ;
        RECT 142.200 94.800 142.600 95.600 ;
        RECT 143.000 94.200 143.300 95.900 ;
        RECT 145.400 94.400 145.800 95.200 ;
        RECT 146.100 94.200 146.400 95.900 ;
        RECT 147.000 95.800 147.400 95.900 ;
        RECT 148.200 95.200 148.600 95.400 ;
        RECT 150.200 95.200 150.500 95.900 ;
        RECT 147.800 94.900 148.600 95.200 ;
        RECT 149.400 94.900 150.600 95.200 ;
        RECT 147.800 94.800 148.200 94.900 ;
        RECT 143.000 93.800 143.400 94.200 ;
        RECT 143.800 93.800 144.200 94.200 ;
        RECT 144.600 94.100 145.000 94.200 ;
        RECT 144.600 93.800 145.400 94.100 ;
        RECT 146.100 93.800 147.400 94.200 ;
        RECT 148.600 93.800 149.000 94.600 ;
        RECT 149.400 94.100 149.700 94.900 ;
        RECT 150.200 94.800 150.600 94.900 ;
        RECT 151.000 94.800 151.500 95.200 ;
        RECT 151.100 94.400 151.500 94.800 ;
        RECT 152.000 94.900 152.300 95.900 ;
        RECT 152.000 94.500 152.500 94.900 ;
        RECT 150.200 94.100 150.600 94.200 ;
        RECT 149.400 93.800 150.600 94.100 ;
        RECT 140.600 91.100 141.000 93.200 ;
        RECT 141.400 93.100 141.800 93.200 ;
        RECT 143.000 93.100 143.300 93.800 ;
        RECT 141.400 92.800 143.300 93.100 ;
        RECT 141.300 92.400 141.700 92.800 ;
        RECT 143.000 92.100 143.300 92.800 ;
        RECT 143.800 93.200 144.100 93.800 ;
        RECT 145.000 93.600 145.400 93.800 ;
        RECT 143.800 92.400 144.200 93.200 ;
        RECT 144.700 93.100 146.500 93.300 ;
        RECT 147.000 93.100 147.300 93.800 ;
        RECT 149.400 93.100 149.700 93.800 ;
        RECT 152.000 93.700 152.300 94.500 ;
        RECT 152.800 94.200 153.100 95.900 ;
        RECT 152.600 93.800 153.100 94.200 ;
        RECT 151.000 93.400 152.300 93.700 ;
        RECT 144.600 93.000 146.600 93.100 ;
        RECT 143.000 91.100 143.400 92.100 ;
        RECT 144.600 91.100 145.000 93.000 ;
        RECT 146.200 91.100 146.600 93.000 ;
        RECT 147.000 91.100 147.400 93.100 ;
        RECT 149.400 91.100 149.800 93.100 ;
        RECT 150.200 92.800 150.600 93.200 ;
        RECT 150.100 92.400 150.500 92.800 ;
        RECT 151.000 91.100 151.400 93.400 ;
        RECT 152.800 93.200 153.100 93.800 ;
        RECT 155.800 95.900 156.500 96.200 ;
        RECT 155.800 95.200 156.100 95.900 ;
        RECT 158.200 95.600 158.600 99.900 ;
        RECT 159.000 95.900 159.400 99.900 ;
        RECT 159.800 96.200 160.200 99.900 ;
        RECT 161.400 96.200 161.800 99.900 ;
        RECT 159.800 95.900 161.800 96.200 ;
        RECT 156.600 95.400 158.600 95.600 ;
        RECT 156.500 95.300 158.600 95.400 ;
        RECT 155.800 94.800 156.200 95.200 ;
        RECT 156.500 95.000 156.900 95.300 ;
        RECT 159.100 95.200 159.400 95.900 ;
        RECT 161.000 95.200 161.400 95.400 ;
        RECT 152.600 92.800 153.100 93.200 ;
        RECT 154.200 93.100 154.600 93.200 ;
        RECT 155.800 93.100 156.100 94.800 ;
        RECT 156.500 93.500 156.800 95.000 ;
        RECT 159.000 94.900 160.200 95.200 ;
        RECT 161.000 94.900 161.800 95.200 ;
        RECT 159.000 94.800 159.400 94.900 ;
        RECT 157.200 94.200 157.600 94.600 ;
        RECT 157.300 93.800 157.800 94.200 ;
        RECT 159.900 94.100 160.200 94.900 ;
        RECT 161.400 94.800 161.800 94.900 ;
        RECT 163.000 95.100 163.400 99.900 ;
        RECT 165.000 96.800 165.400 97.200 ;
        RECT 163.800 95.800 164.200 96.600 ;
        RECT 165.000 96.200 165.300 96.800 ;
        RECT 165.700 96.200 166.100 99.900 ;
        RECT 168.200 96.800 168.600 97.200 ;
        RECT 168.200 96.200 168.500 96.800 ;
        RECT 168.900 96.200 169.300 99.900 ;
        RECT 172.300 97.200 172.700 99.900 ;
        RECT 171.800 96.800 172.700 97.200 ;
        RECT 173.000 96.800 173.400 97.200 ;
        RECT 164.600 95.900 165.300 96.200 ;
        RECT 165.600 95.900 166.100 96.200 ;
        RECT 167.800 95.900 168.500 96.200 ;
        RECT 168.800 95.900 169.300 96.200 ;
        RECT 172.300 96.200 172.700 96.800 ;
        RECT 173.100 96.200 173.400 96.800 ;
        RECT 172.300 95.900 172.800 96.200 ;
        RECT 173.100 96.100 173.800 96.200 ;
        RECT 174.200 96.100 174.600 99.900 ;
        RECT 173.100 95.900 174.600 96.100 ;
        RECT 175.000 96.200 175.400 99.900 ;
        RECT 176.600 96.200 177.000 99.900 ;
        RECT 175.000 95.900 177.000 96.200 ;
        RECT 177.400 97.500 177.800 99.500 ;
        RECT 164.600 95.800 165.000 95.900 ;
        RECT 164.600 95.100 164.900 95.800 ;
        RECT 163.000 94.800 164.900 95.100 ;
        RECT 158.200 93.800 160.200 94.100 ;
        RECT 160.600 93.800 161.000 94.600 ;
        RECT 161.400 94.100 161.800 94.200 ;
        RECT 162.200 94.100 162.600 94.200 ;
        RECT 161.400 93.800 162.600 94.100 ;
        RECT 156.500 93.200 157.700 93.500 ;
        RECT 154.200 92.800 156.200 93.100 ;
        RECT 152.600 91.100 153.000 92.800 ;
        RECT 155.800 91.100 156.200 92.800 ;
        RECT 157.400 92.100 157.700 93.200 ;
        RECT 158.200 93.200 158.500 93.800 ;
        RECT 158.200 92.400 158.600 93.200 ;
        RECT 159.000 92.800 159.400 93.200 ;
        RECT 159.900 93.100 160.200 93.800 ;
        RECT 162.200 93.400 162.600 93.800 ;
        RECT 159.100 92.400 159.500 92.800 ;
        RECT 157.400 91.100 157.800 92.100 ;
        RECT 159.800 91.100 160.200 93.100 ;
        RECT 163.000 93.100 163.400 94.800 ;
        RECT 165.600 94.200 165.900 95.900 ;
        RECT 167.800 95.800 168.200 95.900 ;
        RECT 166.200 94.400 166.600 95.200 ;
        RECT 168.800 94.200 169.100 95.900 ;
        RECT 169.400 94.400 169.800 95.200 ;
        RECT 171.800 94.400 172.200 95.200 ;
        RECT 172.500 94.200 172.800 95.900 ;
        RECT 173.400 95.800 174.600 95.900 ;
        RECT 174.300 95.200 174.600 95.800 ;
        RECT 177.400 95.800 177.700 97.500 ;
        RECT 179.500 96.400 179.900 99.900 ;
        RECT 179.500 96.100 180.300 96.400 ;
        RECT 179.800 95.800 180.300 96.100 ;
        RECT 177.400 95.500 179.300 95.800 ;
        RECT 176.200 95.200 176.600 95.400 ;
        RECT 174.200 94.900 175.400 95.200 ;
        RECT 176.200 94.900 177.000 95.200 ;
        RECT 174.200 94.800 174.600 94.900 ;
        RECT 164.600 93.800 165.900 94.200 ;
        RECT 167.000 94.100 167.400 94.200 ;
        RECT 166.600 93.800 167.400 94.100 ;
        RECT 167.800 93.800 169.100 94.200 ;
        RECT 170.200 94.100 170.600 94.200 ;
        RECT 169.800 93.800 170.600 94.100 ;
        RECT 171.000 94.100 171.400 94.200 ;
        RECT 171.000 93.800 171.800 94.100 ;
        RECT 172.500 93.800 173.800 94.200 ;
        RECT 164.700 93.100 165.000 93.800 ;
        RECT 166.600 93.600 167.000 93.800 ;
        RECT 165.500 93.100 167.300 93.300 ;
        RECT 167.900 93.100 168.200 93.800 ;
        RECT 169.800 93.600 170.200 93.800 ;
        RECT 171.400 93.600 171.800 93.800 ;
        RECT 168.700 93.100 170.500 93.300 ;
        RECT 171.100 93.100 172.900 93.300 ;
        RECT 173.400 93.100 173.700 93.800 ;
        RECT 163.000 92.800 163.900 93.100 ;
        RECT 163.500 91.100 163.900 92.800 ;
        RECT 164.600 91.100 165.000 93.100 ;
        RECT 165.400 93.000 167.400 93.100 ;
        RECT 165.400 91.100 165.800 93.000 ;
        RECT 167.000 91.100 167.400 93.000 ;
        RECT 167.800 91.100 168.200 93.100 ;
        RECT 168.600 93.000 170.600 93.100 ;
        RECT 168.600 91.100 169.000 93.000 ;
        RECT 170.200 91.100 170.600 93.000 ;
        RECT 171.000 93.000 173.000 93.100 ;
        RECT 171.000 91.100 171.400 93.000 ;
        RECT 172.600 91.100 173.000 93.000 ;
        RECT 173.400 91.100 173.800 93.100 ;
        RECT 174.200 92.800 174.600 93.200 ;
        RECT 175.100 93.100 175.400 94.900 ;
        RECT 176.600 94.800 177.000 94.900 ;
        RECT 175.800 93.800 176.200 94.600 ;
        RECT 177.400 94.400 177.800 95.200 ;
        RECT 178.200 94.400 178.600 95.200 ;
        RECT 179.000 94.500 179.300 95.500 ;
        RECT 179.000 94.100 179.700 94.500 ;
        RECT 180.000 94.200 180.300 95.800 ;
        RECT 180.600 94.800 181.000 95.600 ;
        RECT 179.000 93.900 179.500 94.100 ;
        RECT 174.300 92.400 174.700 92.800 ;
        RECT 175.000 91.100 175.400 93.100 ;
        RECT 177.400 93.600 179.500 93.900 ;
        RECT 180.000 93.800 181.000 94.200 ;
        RECT 177.400 92.500 177.700 93.600 ;
        RECT 180.000 93.500 180.300 93.800 ;
        RECT 179.900 93.300 180.300 93.500 ;
        RECT 179.500 93.000 180.300 93.300 ;
        RECT 177.400 91.500 177.800 92.500 ;
        RECT 179.500 91.500 179.900 93.000 ;
        RECT 182.200 91.100 182.600 99.900 ;
        RECT 183.800 95.600 184.200 99.900 ;
        RECT 185.900 97.900 186.500 99.900 ;
        RECT 188.200 97.900 188.600 99.900 ;
        RECT 190.400 98.200 190.800 99.900 ;
        RECT 190.400 97.900 191.400 98.200 ;
        RECT 186.200 97.500 186.600 97.900 ;
        RECT 188.300 97.600 188.600 97.900 ;
        RECT 187.900 97.300 189.700 97.600 ;
        RECT 191.000 97.500 191.400 97.900 ;
        RECT 187.900 97.200 188.300 97.300 ;
        RECT 189.300 97.200 189.700 97.300 ;
        RECT 185.400 97.000 186.100 97.200 ;
        RECT 185.400 96.800 186.500 97.000 ;
        RECT 185.800 96.600 186.500 96.800 ;
        RECT 186.200 96.100 186.500 96.600 ;
        RECT 187.300 96.500 188.400 96.800 ;
        RECT 187.300 96.400 187.700 96.500 ;
        RECT 186.200 95.800 187.400 96.100 ;
        RECT 183.800 95.300 185.900 95.600 ;
        RECT 183.800 93.600 184.200 95.300 ;
        RECT 185.500 95.200 185.900 95.300 ;
        RECT 184.700 94.900 185.100 95.000 ;
        RECT 184.700 94.600 186.600 94.900 ;
        RECT 186.200 94.500 186.600 94.600 ;
        RECT 187.100 94.200 187.400 95.800 ;
        RECT 188.100 95.900 188.400 96.500 ;
        RECT 188.700 96.500 189.100 96.600 ;
        RECT 191.000 96.500 191.400 96.600 ;
        RECT 188.700 96.200 191.400 96.500 ;
        RECT 188.100 95.700 190.500 95.900 ;
        RECT 192.600 95.700 193.000 99.900 ;
        RECT 188.100 95.600 193.000 95.700 ;
        RECT 190.100 95.500 193.000 95.600 ;
        RECT 190.200 95.400 193.000 95.500 ;
        RECT 189.400 95.100 189.800 95.200 ;
        RECT 189.400 94.800 191.900 95.100 ;
        RECT 191.500 94.700 191.900 94.800 ;
        RECT 190.700 94.200 191.100 94.300 ;
        RECT 187.100 93.900 192.600 94.200 ;
        RECT 187.300 93.800 187.700 93.900 ;
        RECT 189.400 93.800 189.800 93.900 ;
        RECT 183.800 93.300 185.700 93.600 ;
        RECT 183.000 93.100 183.400 93.200 ;
        RECT 183.800 93.100 184.200 93.300 ;
        RECT 185.300 93.200 185.700 93.300 ;
        RECT 183.000 92.800 184.200 93.100 ;
        RECT 190.200 92.800 190.500 93.900 ;
        RECT 191.800 93.800 192.600 93.900 ;
        RECT 183.000 92.400 183.400 92.800 ;
        RECT 183.800 91.100 184.200 92.800 ;
        RECT 189.300 92.700 189.700 92.800 ;
        RECT 186.200 92.100 186.600 92.500 ;
        RECT 188.300 92.400 189.700 92.700 ;
        RECT 190.200 92.400 190.600 92.800 ;
        RECT 188.300 92.100 188.600 92.400 ;
        RECT 191.000 92.100 191.400 92.500 ;
        RECT 185.900 91.800 186.600 92.100 ;
        RECT 185.900 91.100 186.500 91.800 ;
        RECT 188.200 91.100 188.600 92.100 ;
        RECT 190.400 91.800 191.400 92.100 ;
        RECT 190.400 91.100 190.800 91.800 ;
        RECT 192.600 91.100 193.000 93.500 ;
        RECT 193.400 91.100 193.800 99.900 ;
        RECT 195.000 95.600 195.400 99.900 ;
        RECT 197.100 97.900 197.700 99.900 ;
        RECT 199.400 97.900 199.800 99.900 ;
        RECT 201.600 98.200 202.000 99.900 ;
        RECT 201.600 97.900 202.600 98.200 ;
        RECT 197.400 97.500 197.800 97.900 ;
        RECT 199.500 97.600 199.800 97.900 ;
        RECT 199.100 97.300 200.900 97.600 ;
        RECT 202.200 97.500 202.600 97.900 ;
        RECT 199.100 97.200 199.500 97.300 ;
        RECT 200.500 97.200 200.900 97.300 ;
        RECT 197.000 96.600 197.700 97.000 ;
        RECT 197.400 96.100 197.700 96.600 ;
        RECT 198.500 96.500 199.600 96.800 ;
        RECT 198.500 96.400 198.900 96.500 ;
        RECT 197.400 95.800 198.600 96.100 ;
        RECT 195.000 95.300 197.100 95.600 ;
        RECT 195.000 93.600 195.400 95.300 ;
        RECT 196.700 95.200 197.100 95.300 ;
        RECT 198.300 95.200 198.600 95.800 ;
        RECT 199.300 95.900 199.600 96.500 ;
        RECT 199.900 96.500 200.300 96.600 ;
        RECT 202.200 96.500 202.600 96.600 ;
        RECT 199.900 96.200 202.600 96.500 ;
        RECT 199.300 95.700 201.700 95.900 ;
        RECT 203.800 95.700 204.200 99.900 ;
        RECT 199.300 95.600 204.200 95.700 ;
        RECT 201.300 95.500 204.200 95.600 ;
        RECT 201.400 95.400 204.200 95.500 ;
        RECT 195.900 94.900 196.300 95.000 ;
        RECT 195.900 94.600 197.800 94.900 ;
        RECT 198.200 94.800 198.600 95.200 ;
        RECT 200.600 95.100 201.000 95.200 ;
        RECT 200.600 94.800 203.100 95.100 ;
        RECT 197.400 94.500 197.800 94.600 ;
        RECT 198.300 94.200 198.600 94.800 ;
        RECT 202.700 94.700 203.100 94.800 ;
        RECT 201.900 94.200 202.300 94.300 ;
        RECT 198.300 93.900 203.800 94.200 ;
        RECT 198.500 93.800 198.900 93.900 ;
        RECT 195.000 93.300 196.900 93.600 ;
        RECT 194.200 93.100 194.600 93.200 ;
        RECT 195.000 93.100 195.400 93.300 ;
        RECT 196.500 93.200 196.900 93.300 ;
        RECT 201.400 93.200 201.700 93.900 ;
        RECT 203.000 93.800 203.800 93.900 ;
        RECT 194.200 92.800 195.400 93.100 ;
        RECT 194.200 92.400 194.600 92.800 ;
        RECT 195.000 91.100 195.400 92.800 ;
        RECT 200.500 92.700 200.900 92.800 ;
        RECT 197.400 92.100 197.800 92.500 ;
        RECT 199.500 92.400 200.900 92.700 ;
        RECT 201.400 92.400 201.800 93.200 ;
        RECT 199.500 92.100 199.800 92.400 ;
        RECT 202.200 92.100 202.600 92.500 ;
        RECT 197.100 91.800 197.800 92.100 ;
        RECT 197.100 91.100 197.700 91.800 ;
        RECT 199.400 91.100 199.800 92.100 ;
        RECT 201.600 91.800 202.600 92.100 ;
        RECT 201.600 91.100 202.000 91.800 ;
        RECT 203.800 91.100 204.200 93.500 ;
        RECT 0.600 87.700 1.000 89.900 ;
        RECT 2.700 89.200 3.300 89.900 ;
        RECT 2.700 88.900 3.400 89.200 ;
        RECT 5.000 88.900 5.400 89.900 ;
        RECT 7.200 89.200 7.600 89.900 ;
        RECT 7.200 88.900 8.200 89.200 ;
        RECT 3.000 88.500 3.400 88.900 ;
        RECT 5.100 88.600 5.400 88.900 ;
        RECT 5.100 88.300 6.500 88.600 ;
        RECT 6.100 88.200 6.500 88.300 ;
        RECT 7.000 88.200 7.400 88.600 ;
        RECT 7.800 88.500 8.200 88.900 ;
        RECT 2.100 87.700 2.500 87.800 ;
        RECT 0.600 87.400 2.500 87.700 ;
        RECT 0.600 85.700 1.000 87.400 ;
        RECT 4.100 87.100 4.500 87.200 ;
        RECT 6.200 87.100 6.600 87.200 ;
        RECT 7.000 87.100 7.300 88.200 ;
        RECT 9.400 87.500 9.800 89.900 ;
        RECT 11.500 88.200 11.900 89.900 ;
        RECT 11.000 87.900 11.900 88.200 ;
        RECT 12.600 87.900 13.000 89.900 ;
        RECT 13.400 88.000 13.800 89.900 ;
        RECT 15.000 88.000 15.400 89.900 ;
        RECT 13.400 87.900 15.400 88.000 ;
        RECT 16.100 88.200 16.500 89.900 ;
        RECT 16.100 87.900 17.000 88.200 ;
        RECT 8.600 87.100 9.400 87.200 ;
        RECT 3.900 86.800 9.400 87.100 ;
        RECT 10.200 86.800 10.600 87.600 ;
        RECT 3.000 86.400 3.400 86.500 ;
        RECT 1.500 86.100 3.400 86.400 ;
        RECT 1.500 86.000 1.900 86.100 ;
        RECT 2.300 85.700 2.700 85.800 ;
        RECT 0.600 85.400 2.700 85.700 ;
        RECT 0.600 81.100 1.000 85.400 ;
        RECT 3.900 85.200 4.200 86.800 ;
        RECT 7.500 86.700 7.900 86.800 ;
        RECT 7.000 86.200 7.400 86.300 ;
        RECT 8.300 86.200 8.700 86.300 ;
        RECT 6.200 85.900 8.700 86.200 ;
        RECT 11.000 86.100 11.400 87.900 ;
        RECT 12.700 87.200 13.000 87.900 ;
        RECT 13.500 87.700 15.300 87.900 ;
        RECT 14.600 87.200 15.000 87.400 ;
        RECT 11.800 87.100 12.200 87.200 ;
        RECT 12.600 87.100 13.900 87.200 ;
        RECT 11.800 86.800 13.900 87.100 ;
        RECT 14.600 87.100 15.400 87.200 ;
        RECT 15.800 87.100 16.200 87.200 ;
        RECT 14.600 86.900 16.200 87.100 ;
        RECT 15.000 86.800 16.200 86.900 ;
        RECT 6.200 85.800 6.600 85.900 ;
        RECT 11.000 85.800 12.900 86.100 ;
        RECT 7.000 85.500 9.800 85.600 ;
        RECT 6.900 85.400 9.800 85.500 ;
        RECT 3.000 84.900 4.200 85.200 ;
        RECT 4.900 85.300 9.800 85.400 ;
        RECT 4.900 85.100 7.300 85.300 ;
        RECT 3.000 84.400 3.300 84.900 ;
        RECT 2.600 84.000 3.300 84.400 ;
        RECT 4.100 84.500 4.500 84.600 ;
        RECT 4.900 84.500 5.200 85.100 ;
        RECT 4.100 84.200 5.200 84.500 ;
        RECT 5.500 84.500 8.200 84.800 ;
        RECT 5.500 84.400 5.900 84.500 ;
        RECT 7.800 84.400 8.200 84.500 ;
        RECT 4.700 83.700 5.100 83.800 ;
        RECT 6.100 83.700 6.500 83.800 ;
        RECT 3.000 83.100 3.400 83.500 ;
        RECT 4.700 83.400 6.500 83.700 ;
        RECT 5.100 83.100 5.400 83.400 ;
        RECT 7.800 83.100 8.200 83.500 ;
        RECT 2.700 81.100 3.300 83.100 ;
        RECT 5.000 81.100 5.400 83.100 ;
        RECT 7.200 82.800 8.200 83.100 ;
        RECT 7.200 81.100 7.600 82.800 ;
        RECT 9.400 81.100 9.800 85.300 ;
        RECT 11.000 81.100 11.400 85.800 ;
        RECT 12.600 85.200 12.900 85.800 ;
        RECT 11.800 84.400 12.200 85.200 ;
        RECT 12.600 85.100 13.000 85.200 ;
        RECT 13.600 85.100 13.900 86.800 ;
        RECT 14.200 85.800 14.600 86.600 ;
        RECT 12.600 84.800 13.300 85.100 ;
        RECT 13.600 84.800 14.100 85.100 ;
        RECT 13.000 84.200 13.300 84.800 ;
        RECT 13.000 83.800 13.400 84.200 ;
        RECT 13.700 81.100 14.100 84.800 ;
        RECT 15.800 84.400 16.200 85.200 ;
        RECT 16.600 81.100 17.000 87.900 ;
        RECT 19.800 87.900 20.200 89.900 ;
        RECT 20.500 88.200 20.900 88.600 ;
        RECT 17.400 86.800 17.800 87.600 ;
        RECT 19.000 86.400 19.400 87.200 ;
        RECT 18.200 86.100 18.600 86.200 ;
        RECT 19.800 86.100 20.100 87.900 ;
        RECT 20.600 87.800 21.000 88.200 ;
        RECT 21.400 87.900 21.800 89.900 ;
        RECT 22.200 88.000 22.600 89.900 ;
        RECT 23.800 88.000 24.200 89.900 ;
        RECT 22.200 87.900 24.200 88.000 ;
        RECT 21.500 87.200 21.800 87.900 ;
        RECT 22.300 87.700 24.100 87.900 ;
        RECT 24.600 87.500 25.000 89.900 ;
        RECT 26.800 89.200 27.200 89.900 ;
        RECT 26.200 88.900 27.200 89.200 ;
        RECT 29.000 88.900 29.400 89.900 ;
        RECT 31.100 89.200 31.700 89.900 ;
        RECT 31.000 88.900 31.700 89.200 ;
        RECT 26.200 88.500 26.600 88.900 ;
        RECT 29.000 88.600 29.300 88.900 ;
        RECT 27.000 88.200 27.400 88.600 ;
        RECT 27.900 88.300 29.300 88.600 ;
        RECT 31.000 88.500 31.400 88.900 ;
        RECT 27.900 88.200 28.300 88.300 ;
        RECT 23.400 87.200 23.800 87.400 ;
        RECT 21.400 86.800 22.700 87.200 ;
        RECT 23.400 86.900 24.200 87.200 ;
        RECT 23.800 86.800 24.200 86.900 ;
        RECT 25.000 87.100 25.800 87.200 ;
        RECT 27.100 87.100 27.400 88.200 ;
        RECT 33.400 88.100 33.800 89.900 ;
        RECT 35.000 88.900 35.400 89.900 ;
        RECT 34.200 88.100 34.600 88.600 ;
        RECT 35.100 88.100 35.400 88.900 ;
        RECT 36.700 88.200 37.100 88.600 ;
        RECT 36.600 88.100 37.000 88.200 ;
        RECT 33.400 87.800 34.600 88.100 ;
        RECT 35.000 87.800 37.000 88.100 ;
        RECT 37.400 87.800 37.800 89.900 ;
        RECT 31.900 87.700 32.300 87.800 ;
        RECT 33.400 87.700 33.800 87.800 ;
        RECT 31.900 87.400 33.800 87.700 ;
        RECT 29.400 87.100 30.300 87.200 ;
        RECT 25.000 86.800 30.500 87.100 ;
        RECT 20.600 86.100 21.000 86.200 ;
        RECT 18.200 85.800 19.000 86.100 ;
        RECT 19.800 85.800 21.000 86.100 ;
        RECT 18.600 85.600 19.000 85.800 ;
        RECT 20.600 85.100 20.900 85.800 ;
        RECT 21.400 85.100 21.800 85.200 ;
        RECT 22.400 85.100 22.700 86.800 ;
        RECT 26.500 86.700 26.900 86.800 ;
        RECT 23.000 85.800 23.400 86.600 ;
        RECT 25.700 86.200 26.100 86.300 ;
        RECT 25.700 85.900 28.200 86.200 ;
        RECT 27.800 85.800 28.200 85.900 ;
        RECT 24.600 85.500 27.400 85.600 ;
        RECT 24.600 85.400 27.500 85.500 ;
        RECT 24.600 85.300 29.500 85.400 ;
        RECT 18.200 84.800 20.200 85.100 ;
        RECT 18.200 81.100 18.600 84.800 ;
        RECT 19.800 81.100 20.200 84.800 ;
        RECT 20.600 84.800 22.100 85.100 ;
        RECT 22.400 84.800 22.900 85.100 ;
        RECT 20.600 81.100 21.000 84.800 ;
        RECT 21.800 84.200 22.100 84.800 ;
        RECT 21.800 83.800 22.200 84.200 ;
        RECT 22.500 81.100 22.900 84.800 ;
        RECT 24.600 81.100 25.000 85.300 ;
        RECT 27.100 85.100 29.500 85.300 ;
        RECT 26.200 84.500 28.900 84.800 ;
        RECT 26.200 84.400 26.600 84.500 ;
        RECT 28.500 84.400 28.900 84.500 ;
        RECT 29.200 84.500 29.500 85.100 ;
        RECT 30.200 85.200 30.500 86.800 ;
        RECT 31.000 86.400 31.400 86.500 ;
        RECT 31.000 86.100 32.900 86.400 ;
        RECT 32.500 86.000 32.900 86.100 ;
        RECT 33.400 86.100 33.800 87.400 ;
        RECT 35.100 87.200 35.400 87.800 ;
        RECT 34.200 86.800 34.600 87.200 ;
        RECT 35.000 86.800 35.400 87.200 ;
        RECT 34.200 86.100 34.500 86.800 ;
        RECT 33.400 85.800 34.500 86.100 ;
        RECT 31.700 85.700 32.100 85.800 ;
        RECT 33.400 85.700 33.800 85.800 ;
        RECT 31.700 85.400 33.800 85.700 ;
        RECT 30.200 84.900 31.400 85.200 ;
        RECT 29.900 84.500 30.300 84.600 ;
        RECT 29.200 84.200 30.300 84.500 ;
        RECT 31.100 84.400 31.400 84.900 ;
        RECT 31.100 84.000 31.800 84.400 ;
        RECT 27.900 83.700 28.300 83.800 ;
        RECT 29.300 83.700 29.700 83.800 ;
        RECT 26.200 83.100 26.600 83.500 ;
        RECT 27.900 83.400 29.700 83.700 ;
        RECT 29.000 83.100 29.300 83.400 ;
        RECT 31.000 83.100 31.400 83.500 ;
        RECT 26.200 82.800 27.200 83.100 ;
        RECT 26.800 81.100 27.200 82.800 ;
        RECT 29.000 81.100 29.400 83.100 ;
        RECT 31.100 81.100 31.700 83.100 ;
        RECT 33.400 81.100 33.800 85.400 ;
        RECT 35.100 85.100 35.400 86.800 ;
        RECT 35.800 85.400 36.200 86.200 ;
        RECT 36.600 86.100 37.000 86.200 ;
        RECT 37.500 86.100 37.800 87.800 ;
        RECT 41.400 87.900 41.800 89.900 ;
        RECT 42.100 88.200 42.500 88.600 ;
        RECT 38.200 86.400 38.600 87.200 ;
        RECT 40.600 86.400 41.000 87.200 ;
        RECT 39.000 86.100 39.400 86.200 ;
        RECT 36.600 85.800 37.800 86.100 ;
        RECT 38.600 85.800 39.400 86.100 ;
        RECT 39.800 86.100 40.200 86.200 ;
        RECT 41.400 86.100 41.700 87.900 ;
        RECT 42.200 87.800 42.600 88.200 ;
        RECT 43.000 87.900 43.400 89.900 ;
        RECT 43.800 88.000 44.200 89.900 ;
        RECT 45.400 88.000 45.800 89.900 ;
        RECT 43.800 87.900 45.800 88.000 ;
        RECT 43.100 87.200 43.400 87.900 ;
        RECT 43.900 87.700 45.700 87.900 ;
        RECT 45.000 87.200 45.400 87.400 ;
        RECT 43.000 86.800 44.300 87.200 ;
        RECT 45.000 86.900 45.800 87.200 ;
        RECT 45.400 86.800 45.800 86.900 ;
        RECT 42.200 86.100 42.600 86.200 ;
        RECT 39.800 85.800 40.600 86.100 ;
        RECT 41.400 85.800 42.600 86.100 ;
        RECT 36.700 85.100 37.000 85.800 ;
        RECT 38.600 85.600 39.000 85.800 ;
        RECT 40.200 85.600 40.600 85.800 ;
        RECT 42.200 85.100 42.500 85.800 ;
        RECT 43.000 85.100 43.400 85.200 ;
        RECT 44.000 85.100 44.300 86.800 ;
        RECT 44.600 86.100 45.000 86.600 ;
        RECT 46.200 86.100 46.600 89.900 ;
        RECT 47.000 88.100 47.400 88.600 ;
        RECT 49.400 88.100 49.800 89.900 ;
        RECT 51.500 89.200 52.100 89.900 ;
        RECT 51.500 88.900 52.200 89.200 ;
        RECT 53.800 88.900 54.200 89.900 ;
        RECT 56.000 89.200 56.400 89.900 ;
        RECT 56.000 88.900 57.000 89.200 ;
        RECT 51.800 88.500 52.200 88.900 ;
        RECT 53.900 88.600 54.200 88.900 ;
        RECT 53.900 88.300 55.300 88.600 ;
        RECT 54.900 88.200 55.300 88.300 ;
        RECT 47.000 87.800 49.800 88.100 ;
        RECT 55.800 87.800 56.200 88.600 ;
        RECT 56.600 88.500 57.000 88.900 ;
        RECT 44.600 85.800 46.600 86.100 ;
        RECT 35.000 84.700 35.900 85.100 ;
        RECT 35.500 81.100 35.900 84.700 ;
        RECT 36.600 81.100 37.000 85.100 ;
        RECT 37.400 84.800 39.400 85.100 ;
        RECT 37.400 81.100 37.800 84.800 ;
        RECT 39.000 81.100 39.400 84.800 ;
        RECT 39.800 84.800 41.800 85.100 ;
        RECT 39.800 81.100 40.200 84.800 ;
        RECT 41.400 81.100 41.800 84.800 ;
        RECT 42.200 84.800 43.700 85.100 ;
        RECT 44.000 84.800 44.500 85.100 ;
        RECT 42.200 81.100 42.600 84.800 ;
        RECT 43.400 84.200 43.700 84.800 ;
        RECT 43.400 83.800 43.800 84.200 ;
        RECT 44.100 81.100 44.500 84.800 ;
        RECT 46.200 81.100 46.600 85.800 ;
        RECT 49.400 87.700 49.800 87.800 ;
        RECT 50.900 87.700 51.300 87.800 ;
        RECT 49.400 87.400 51.300 87.700 ;
        RECT 49.400 85.700 49.800 87.400 ;
        RECT 52.900 87.100 53.300 87.200 ;
        RECT 55.800 87.100 56.100 87.800 ;
        RECT 58.200 87.500 58.600 89.900 ;
        RECT 60.300 88.200 60.700 89.900 ;
        RECT 59.800 87.900 60.700 88.200 ;
        RECT 61.400 87.900 61.800 89.900 ;
        RECT 62.200 88.000 62.600 89.900 ;
        RECT 63.800 88.000 64.200 89.900 ;
        RECT 62.200 87.900 64.200 88.000 ;
        RECT 57.400 87.100 58.200 87.200 ;
        RECT 52.700 86.800 58.200 87.100 ;
        RECT 59.000 86.800 59.400 87.600 ;
        RECT 51.800 86.400 52.200 86.500 ;
        RECT 50.300 86.100 52.200 86.400 ;
        RECT 50.300 86.000 50.700 86.100 ;
        RECT 51.100 85.700 51.500 85.800 ;
        RECT 49.400 85.400 51.500 85.700 ;
        RECT 49.400 81.100 49.800 85.400 ;
        RECT 52.700 85.200 53.000 86.800 ;
        RECT 56.300 86.700 56.700 86.800 ;
        RECT 55.800 86.200 56.200 86.300 ;
        RECT 57.100 86.200 57.500 86.300 ;
        RECT 55.000 85.900 57.500 86.200 ;
        RECT 59.800 86.100 60.200 87.900 ;
        RECT 61.500 87.200 61.800 87.900 ;
        RECT 62.300 87.700 64.100 87.900 ;
        RECT 64.600 87.600 65.000 89.900 ;
        RECT 66.200 88.200 66.600 89.900 ;
        RECT 66.200 87.900 66.700 88.200 ;
        RECT 67.800 87.900 68.200 89.900 ;
        RECT 68.600 88.000 69.000 89.900 ;
        RECT 70.200 88.000 70.600 89.900 ;
        RECT 68.600 87.900 70.600 88.000 ;
        RECT 71.000 87.900 71.400 89.900 ;
        RECT 71.800 88.000 72.200 89.900 ;
        RECT 73.400 88.000 73.800 89.900 ;
        RECT 74.300 88.200 74.700 88.600 ;
        RECT 71.800 87.900 73.800 88.000 ;
        RECT 63.400 87.200 63.800 87.400 ;
        RECT 64.600 87.300 65.900 87.600 ;
        RECT 60.600 87.100 61.000 87.200 ;
        RECT 61.400 87.100 62.700 87.200 ;
        RECT 60.600 86.800 62.700 87.100 ;
        RECT 63.400 86.900 64.200 87.200 ;
        RECT 63.800 86.800 64.200 86.900 ;
        RECT 55.000 85.800 55.400 85.900 ;
        RECT 59.800 85.800 61.700 86.100 ;
        RECT 55.800 85.500 58.600 85.600 ;
        RECT 55.700 85.400 58.600 85.500 ;
        RECT 51.800 84.900 53.000 85.200 ;
        RECT 53.700 85.300 58.600 85.400 ;
        RECT 53.700 85.100 56.100 85.300 ;
        RECT 51.800 84.400 52.100 84.900 ;
        RECT 51.400 84.000 52.100 84.400 ;
        RECT 52.900 84.500 53.300 84.600 ;
        RECT 53.700 84.500 54.000 85.100 ;
        RECT 52.900 84.200 54.000 84.500 ;
        RECT 54.300 84.500 57.000 84.800 ;
        RECT 54.300 84.400 54.700 84.500 ;
        RECT 56.600 84.400 57.000 84.500 ;
        RECT 53.500 83.700 53.900 83.800 ;
        RECT 54.900 83.700 55.300 83.800 ;
        RECT 51.800 83.100 52.200 83.500 ;
        RECT 53.500 83.400 55.300 83.700 ;
        RECT 53.900 83.100 54.200 83.400 ;
        RECT 56.600 83.100 57.000 83.500 ;
        RECT 51.500 81.100 52.100 83.100 ;
        RECT 53.800 81.100 54.200 83.100 ;
        RECT 56.000 82.800 57.000 83.100 ;
        RECT 56.000 81.100 56.400 82.800 ;
        RECT 58.200 81.100 58.600 85.300 ;
        RECT 59.800 81.100 60.200 85.800 ;
        RECT 61.400 85.200 61.700 85.800 ;
        RECT 60.600 84.400 61.000 85.200 ;
        RECT 61.400 85.100 61.800 85.200 ;
        RECT 62.400 85.100 62.700 86.800 ;
        RECT 63.000 85.800 63.400 86.600 ;
        RECT 64.700 86.200 65.100 86.600 ;
        RECT 64.600 85.800 65.100 86.200 ;
        RECT 65.600 86.500 65.900 87.300 ;
        RECT 66.400 87.200 66.700 87.900 ;
        RECT 67.900 87.200 68.200 87.900 ;
        RECT 68.700 87.700 70.500 87.900 ;
        RECT 69.800 87.200 70.200 87.400 ;
        RECT 71.100 87.200 71.400 87.900 ;
        RECT 71.900 87.700 73.700 87.900 ;
        RECT 74.200 87.800 74.600 88.200 ;
        RECT 75.000 87.900 75.400 89.900 ;
        RECT 78.200 88.200 78.600 89.900 ;
        RECT 73.000 87.200 73.400 87.400 ;
        RECT 66.200 86.800 66.700 87.200 ;
        RECT 67.800 86.800 69.100 87.200 ;
        RECT 69.800 86.900 70.600 87.200 ;
        RECT 70.200 86.800 70.600 86.900 ;
        RECT 71.000 86.800 72.300 87.200 ;
        RECT 73.000 86.900 73.800 87.200 ;
        RECT 73.400 86.800 73.800 86.900 ;
        RECT 65.600 86.100 66.100 86.500 ;
        RECT 65.600 85.100 65.900 86.100 ;
        RECT 66.400 85.100 66.700 86.800 ;
        RECT 67.000 86.100 67.400 86.200 ;
        RECT 67.000 85.800 68.100 86.100 ;
        RECT 61.400 84.800 62.100 85.100 ;
        RECT 62.400 84.800 62.900 85.100 ;
        RECT 61.800 84.200 62.100 84.800 ;
        RECT 61.800 83.800 62.200 84.200 ;
        RECT 62.500 81.100 62.900 84.800 ;
        RECT 64.600 84.800 65.900 85.100 ;
        RECT 64.600 81.100 65.000 84.800 ;
        RECT 66.200 84.600 66.700 85.100 ;
        RECT 67.800 85.200 68.100 85.800 ;
        RECT 67.800 85.100 68.200 85.200 ;
        RECT 68.800 85.100 69.100 86.800 ;
        RECT 69.400 85.800 69.800 86.600 ;
        RECT 71.000 85.100 71.400 85.200 ;
        RECT 72.000 85.100 72.300 86.800 ;
        RECT 72.600 86.100 73.000 86.600 ;
        RECT 73.400 86.100 73.800 86.200 ;
        RECT 72.600 85.800 73.800 86.100 ;
        RECT 74.200 86.100 74.600 86.200 ;
        RECT 75.100 86.100 75.400 87.900 ;
        RECT 78.100 87.900 78.600 88.200 ;
        RECT 78.100 87.200 78.400 87.900 ;
        RECT 79.800 87.600 80.200 89.900 ;
        RECT 80.600 88.000 81.000 89.900 ;
        RECT 82.200 88.000 82.600 89.900 ;
        RECT 80.600 87.900 82.600 88.000 ;
        RECT 83.000 87.900 83.400 89.900 ;
        RECT 83.800 87.900 84.200 89.900 ;
        RECT 84.600 88.000 85.000 89.900 ;
        RECT 86.200 88.000 86.600 89.900 ;
        RECT 84.600 87.900 86.600 88.000 ;
        RECT 80.700 87.700 82.500 87.900 ;
        RECT 78.900 87.300 80.200 87.600 ;
        RECT 75.800 86.400 76.200 87.200 ;
        RECT 78.100 86.800 78.600 87.200 ;
        RECT 76.600 86.100 77.000 86.200 ;
        RECT 74.200 85.800 75.400 86.100 ;
        RECT 76.200 85.800 77.000 86.100 ;
        RECT 74.300 85.100 74.600 85.800 ;
        RECT 76.200 85.600 76.600 85.800 ;
        RECT 78.100 85.200 78.400 86.800 ;
        RECT 78.900 86.500 79.200 87.300 ;
        RECT 81.000 87.200 81.400 87.400 ;
        RECT 83.000 87.200 83.300 87.900 ;
        RECT 83.900 87.200 84.200 87.900 ;
        RECT 84.700 87.700 86.500 87.900 ;
        RECT 87.800 87.600 88.200 89.900 ;
        RECT 89.400 87.600 89.800 89.900 ;
        RECT 85.800 87.200 86.200 87.400 ;
        RECT 80.600 86.900 81.400 87.200 ;
        RECT 80.600 86.800 81.000 86.900 ;
        RECT 82.100 86.800 83.400 87.200 ;
        RECT 83.800 86.800 85.100 87.200 ;
        RECT 85.800 86.900 86.600 87.200 ;
        RECT 86.200 86.800 86.600 86.900 ;
        RECT 87.000 86.800 87.400 87.600 ;
        RECT 87.800 87.200 89.800 87.600 ;
        RECT 92.600 87.900 93.000 89.900 ;
        RECT 93.300 88.200 93.700 88.600 ;
        RECT 78.700 86.100 79.200 86.500 ;
        RECT 67.800 84.800 68.500 85.100 ;
        RECT 68.800 84.800 69.300 85.100 ;
        RECT 71.000 84.800 71.700 85.100 ;
        RECT 72.000 84.800 72.500 85.100 ;
        RECT 66.200 81.100 66.600 84.600 ;
        RECT 68.200 84.200 68.500 84.800 ;
        RECT 67.800 83.800 68.600 84.200 ;
        RECT 68.900 81.100 69.300 84.800 ;
        RECT 71.400 84.200 71.700 84.800 ;
        RECT 71.400 83.800 71.800 84.200 ;
        RECT 72.100 83.200 72.500 84.800 ;
        RECT 72.100 82.800 73.000 83.200 ;
        RECT 72.100 81.100 72.500 82.800 ;
        RECT 74.200 81.100 74.600 85.100 ;
        RECT 75.000 84.800 77.000 85.100 ;
        RECT 75.000 81.100 75.400 84.800 ;
        RECT 76.600 81.100 77.000 84.800 ;
        RECT 78.100 84.600 78.600 85.200 ;
        RECT 78.900 85.100 79.200 86.100 ;
        RECT 79.700 86.200 80.100 86.600 ;
        RECT 79.700 85.800 80.200 86.200 ;
        RECT 80.600 86.100 81.000 86.200 ;
        RECT 81.400 86.100 81.800 86.600 ;
        RECT 80.600 85.800 81.800 86.100 ;
        RECT 82.100 85.100 82.400 86.800 ;
        RECT 83.000 85.100 83.400 85.200 ;
        RECT 78.900 84.800 80.200 85.100 ;
        RECT 78.200 81.100 78.600 84.600 ;
        RECT 79.800 81.100 80.200 84.800 ;
        RECT 81.900 84.800 82.400 85.100 ;
        RECT 82.700 84.800 83.400 85.100 ;
        RECT 83.800 85.100 84.200 85.200 ;
        RECT 84.800 85.100 85.100 86.800 ;
        RECT 85.400 85.800 85.800 86.600 ;
        RECT 87.000 86.100 87.400 86.200 ;
        RECT 87.000 85.800 88.200 86.100 ;
        RECT 89.400 85.800 89.800 87.200 ;
        RECT 91.800 86.400 92.200 87.200 ;
        RECT 91.000 86.100 91.400 86.200 ;
        RECT 92.600 86.100 92.900 87.900 ;
        RECT 93.400 87.800 93.800 88.200 ;
        RECT 94.200 87.900 94.600 89.900 ;
        RECT 95.000 88.000 95.400 89.900 ;
        RECT 96.600 88.000 97.000 89.900 ;
        RECT 95.000 87.900 97.000 88.000 ;
        RECT 94.300 87.200 94.600 87.900 ;
        RECT 95.100 87.700 96.900 87.900 ;
        RECT 96.200 87.200 96.600 87.400 ;
        RECT 94.200 86.800 95.500 87.200 ;
        RECT 96.200 86.900 97.000 87.200 ;
        RECT 96.600 86.800 97.000 86.900 ;
        RECT 93.400 86.100 93.800 86.200 ;
        RECT 91.000 85.800 91.800 86.100 ;
        RECT 92.600 85.800 93.800 86.100 ;
        RECT 87.800 85.400 89.800 85.800 ;
        RECT 91.400 85.600 91.800 85.800 ;
        RECT 83.800 84.800 84.500 85.100 ;
        RECT 84.800 84.800 85.300 85.100 ;
        RECT 81.900 81.100 82.300 84.800 ;
        RECT 82.700 84.200 83.000 84.800 ;
        RECT 82.600 83.800 83.000 84.200 ;
        RECT 84.200 84.200 84.500 84.800 ;
        RECT 84.200 83.800 84.600 84.200 ;
        RECT 84.900 81.100 85.300 84.800 ;
        RECT 87.800 81.100 88.200 85.400 ;
        RECT 89.400 81.100 89.800 85.400 ;
        RECT 93.400 85.100 93.700 85.800 ;
        RECT 94.200 85.100 94.600 85.200 ;
        RECT 95.200 85.100 95.500 86.800 ;
        RECT 95.800 86.100 96.200 86.600 ;
        RECT 97.400 86.100 97.800 89.900 ;
        RECT 98.200 87.800 98.600 88.600 ;
        RECT 100.300 88.200 100.700 89.900 ;
        RECT 99.800 87.900 100.700 88.200 ;
        RECT 103.000 87.900 103.400 89.900 ;
        RECT 103.800 88.000 104.200 89.900 ;
        RECT 105.400 88.000 105.800 89.900 ;
        RECT 103.800 87.900 105.800 88.000 ;
        RECT 99.000 86.800 99.400 87.600 ;
        RECT 95.800 85.800 97.800 86.100 ;
        RECT 91.000 84.800 93.000 85.100 ;
        RECT 91.000 81.100 91.400 84.800 ;
        RECT 92.600 81.100 93.000 84.800 ;
        RECT 93.400 81.100 93.800 85.100 ;
        RECT 94.200 84.800 94.900 85.100 ;
        RECT 95.200 84.800 95.700 85.100 ;
        RECT 94.600 84.200 94.900 84.800 ;
        RECT 94.600 83.800 95.000 84.200 ;
        RECT 95.300 82.200 95.700 84.800 ;
        RECT 95.300 81.800 96.200 82.200 ;
        RECT 95.300 81.100 95.700 81.800 ;
        RECT 97.400 81.100 97.800 85.800 ;
        RECT 99.800 86.100 100.200 87.900 ;
        RECT 103.100 87.200 103.400 87.900 ;
        RECT 103.900 87.700 105.700 87.900 ;
        RECT 106.200 87.700 106.600 89.900 ;
        RECT 108.300 89.200 108.900 89.900 ;
        RECT 108.300 88.900 109.000 89.200 ;
        RECT 110.600 88.900 111.000 89.900 ;
        RECT 112.800 89.200 113.200 89.900 ;
        RECT 112.800 88.900 113.800 89.200 ;
        RECT 108.600 88.500 109.000 88.900 ;
        RECT 110.700 88.600 111.000 88.900 ;
        RECT 110.700 88.300 112.100 88.600 ;
        RECT 111.700 88.200 112.100 88.300 ;
        RECT 112.600 88.200 113.000 88.600 ;
        RECT 113.400 88.500 113.800 88.900 ;
        RECT 107.700 87.700 108.100 87.800 ;
        RECT 106.200 87.400 108.100 87.700 ;
        RECT 105.000 87.200 105.400 87.400 ;
        RECT 103.000 86.800 104.300 87.200 ;
        RECT 105.000 86.900 105.800 87.200 ;
        RECT 105.400 86.800 105.800 86.900 ;
        RECT 99.800 85.800 103.300 86.100 ;
        RECT 99.800 81.100 100.200 85.800 ;
        RECT 103.000 85.200 103.300 85.800 ;
        RECT 100.600 84.400 101.000 85.200 ;
        RECT 103.000 85.100 103.400 85.200 ;
        RECT 104.000 85.100 104.300 86.800 ;
        RECT 104.600 85.800 105.000 86.600 ;
        RECT 106.200 85.700 106.600 87.400 ;
        RECT 109.700 87.100 110.600 87.200 ;
        RECT 112.600 87.100 112.900 88.200 ;
        RECT 115.000 87.500 115.400 89.900 ;
        RECT 115.900 88.200 116.300 88.600 ;
        RECT 115.800 87.800 116.200 88.200 ;
        RECT 116.600 87.900 117.000 89.900 ;
        RECT 114.200 87.100 115.000 87.200 ;
        RECT 109.500 86.800 115.000 87.100 ;
        RECT 108.600 86.400 109.000 86.500 ;
        RECT 107.100 86.100 109.000 86.400 ;
        RECT 107.100 86.000 107.500 86.100 ;
        RECT 107.900 85.700 108.300 85.800 ;
        RECT 106.200 85.400 108.300 85.700 ;
        RECT 103.000 84.800 103.700 85.100 ;
        RECT 104.000 84.800 104.500 85.100 ;
        RECT 103.400 84.200 103.700 84.800 ;
        RECT 103.400 83.800 103.800 84.200 ;
        RECT 104.100 81.100 104.500 84.800 ;
        RECT 106.200 81.100 106.600 85.400 ;
        RECT 109.500 85.200 109.800 86.800 ;
        RECT 113.100 86.700 113.500 86.800 ;
        RECT 113.900 86.200 114.300 86.300 ;
        RECT 116.700 86.200 117.000 87.900 ;
        RECT 119.000 87.700 119.400 89.900 ;
        RECT 121.100 89.200 121.700 89.900 ;
        RECT 121.100 88.900 121.800 89.200 ;
        RECT 123.400 88.900 123.800 89.900 ;
        RECT 125.600 89.200 126.000 89.900 ;
        RECT 125.600 88.900 126.600 89.200 ;
        RECT 121.400 88.500 121.800 88.900 ;
        RECT 123.500 88.600 123.800 88.900 ;
        RECT 123.500 88.300 124.900 88.600 ;
        RECT 124.500 88.200 124.900 88.300 ;
        RECT 125.400 88.200 125.800 88.600 ;
        RECT 126.200 88.500 126.600 88.900 ;
        RECT 120.500 87.700 120.900 87.800 ;
        RECT 119.000 87.400 120.900 87.700 ;
        RECT 117.400 86.400 117.800 87.200 ;
        RECT 110.200 86.100 110.600 86.200 ;
        RECT 111.800 86.100 114.300 86.200 ;
        RECT 110.200 85.900 114.300 86.100 ;
        RECT 115.800 86.100 116.200 86.200 ;
        RECT 116.600 86.100 117.000 86.200 ;
        RECT 118.200 86.100 118.600 86.200 ;
        RECT 110.200 85.800 112.200 85.900 ;
        RECT 115.800 85.800 117.000 86.100 ;
        RECT 117.800 85.800 118.600 86.100 ;
        RECT 112.600 85.500 115.400 85.600 ;
        RECT 112.500 85.400 115.400 85.500 ;
        RECT 108.600 84.900 109.800 85.200 ;
        RECT 110.500 85.300 115.400 85.400 ;
        RECT 110.500 85.100 112.900 85.300 ;
        RECT 108.600 84.400 108.900 84.900 ;
        RECT 108.200 84.000 108.900 84.400 ;
        RECT 109.700 84.500 110.100 84.600 ;
        RECT 110.500 84.500 110.800 85.100 ;
        RECT 109.700 84.200 110.800 84.500 ;
        RECT 111.100 84.500 113.800 84.800 ;
        RECT 111.100 84.400 111.500 84.500 ;
        RECT 113.400 84.400 113.800 84.500 ;
        RECT 110.300 83.700 110.700 83.800 ;
        RECT 111.700 83.700 112.100 83.800 ;
        RECT 108.600 83.100 109.000 83.500 ;
        RECT 110.300 83.400 112.100 83.700 ;
        RECT 110.700 83.100 111.000 83.400 ;
        RECT 113.400 83.100 113.800 83.500 ;
        RECT 108.300 81.100 108.900 83.100 ;
        RECT 110.600 81.100 111.000 83.100 ;
        RECT 112.800 82.800 113.800 83.100 ;
        RECT 112.800 81.100 113.200 82.800 ;
        RECT 115.000 81.100 115.400 85.300 ;
        RECT 115.900 85.100 116.200 85.800 ;
        RECT 117.800 85.600 118.200 85.800 ;
        RECT 119.000 85.700 119.400 87.400 ;
        RECT 122.500 87.100 122.900 87.200 ;
        RECT 125.400 87.100 125.700 88.200 ;
        RECT 127.800 87.500 128.200 89.900 ;
        RECT 129.400 88.900 129.800 89.900 ;
        RECT 128.600 87.800 129.000 88.600 ;
        RECT 129.500 88.100 129.800 88.900 ;
        RECT 131.100 88.200 131.500 88.600 ;
        RECT 131.000 88.100 131.400 88.200 ;
        RECT 129.400 87.800 131.400 88.100 ;
        RECT 131.800 87.900 132.200 89.900 ;
        RECT 129.500 87.200 129.800 87.800 ;
        RECT 127.000 87.100 127.800 87.200 ;
        RECT 122.300 86.800 127.800 87.100 ;
        RECT 129.400 86.800 129.800 87.200 ;
        RECT 131.000 87.100 131.400 87.200 ;
        RECT 131.900 87.100 132.200 87.900 ;
        RECT 134.200 87.600 134.600 89.900 ;
        RECT 135.800 88.200 136.200 89.900 ;
        RECT 135.800 87.900 136.300 88.200 ;
        RECT 134.200 87.300 135.500 87.600 ;
        RECT 131.000 86.800 132.200 87.100 ;
        RECT 121.400 86.400 121.800 86.500 ;
        RECT 119.900 86.100 121.800 86.400 ;
        RECT 122.300 86.200 122.600 86.800 ;
        RECT 125.900 86.700 126.300 86.800 ;
        RECT 125.400 86.200 125.800 86.300 ;
        RECT 126.700 86.200 127.100 86.300 ;
        RECT 119.900 86.000 120.300 86.100 ;
        RECT 122.200 85.800 122.600 86.200 ;
        RECT 124.600 85.900 127.100 86.200 ;
        RECT 124.600 85.800 125.000 85.900 ;
        RECT 120.700 85.700 121.100 85.800 ;
        RECT 119.000 85.400 121.100 85.700 ;
        RECT 115.800 81.100 116.200 85.100 ;
        RECT 116.600 84.800 118.600 85.100 ;
        RECT 116.600 81.100 117.000 84.800 ;
        RECT 118.200 81.100 118.600 84.800 ;
        RECT 119.000 81.100 119.400 85.400 ;
        RECT 122.300 85.200 122.600 85.800 ;
        RECT 125.400 85.500 128.200 85.600 ;
        RECT 125.300 85.400 128.200 85.500 ;
        RECT 121.400 84.900 122.600 85.200 ;
        RECT 123.300 85.300 128.200 85.400 ;
        RECT 123.300 85.100 125.700 85.300 ;
        RECT 121.400 84.400 121.700 84.900 ;
        RECT 121.000 84.000 121.700 84.400 ;
        RECT 122.500 84.500 122.900 84.600 ;
        RECT 123.300 84.500 123.600 85.100 ;
        RECT 122.500 84.200 123.600 84.500 ;
        RECT 123.900 84.500 126.600 84.800 ;
        RECT 123.900 84.400 124.300 84.500 ;
        RECT 126.200 84.400 126.600 84.500 ;
        RECT 123.100 83.700 123.500 83.800 ;
        RECT 124.500 83.700 124.900 83.800 ;
        RECT 121.400 83.100 121.800 83.500 ;
        RECT 123.100 83.400 124.900 83.700 ;
        RECT 123.500 83.100 123.800 83.400 ;
        RECT 126.200 83.100 126.600 83.500 ;
        RECT 121.100 81.100 121.700 83.100 ;
        RECT 123.400 81.100 123.800 83.100 ;
        RECT 125.600 82.800 126.600 83.100 ;
        RECT 125.600 81.100 126.000 82.800 ;
        RECT 127.800 81.100 128.200 85.300 ;
        RECT 129.500 85.100 129.800 86.800 ;
        RECT 130.200 85.400 130.600 86.200 ;
        RECT 131.000 86.100 131.400 86.200 ;
        RECT 131.900 86.100 132.200 86.800 ;
        RECT 132.600 87.100 133.000 87.200 ;
        RECT 133.400 87.100 133.800 87.200 ;
        RECT 132.600 86.800 133.800 87.100 ;
        RECT 132.600 86.400 133.000 86.800 ;
        RECT 134.300 86.200 134.700 86.600 ;
        RECT 133.400 86.100 133.800 86.200 ;
        RECT 131.000 85.800 132.200 86.100 ;
        RECT 133.000 85.800 133.800 86.100 ;
        RECT 134.200 85.800 134.700 86.200 ;
        RECT 135.200 86.500 135.500 87.300 ;
        RECT 136.000 87.200 136.300 87.900 ;
        RECT 135.800 86.800 136.300 87.200 ;
        RECT 135.200 86.100 135.700 86.500 ;
        RECT 131.100 85.100 131.400 85.800 ;
        RECT 133.000 85.600 133.400 85.800 ;
        RECT 135.200 85.100 135.500 86.100 ;
        RECT 136.000 85.100 136.300 86.800 ;
        RECT 129.400 84.700 130.300 85.100 ;
        RECT 129.900 81.100 130.300 84.700 ;
        RECT 131.000 81.100 131.400 85.100 ;
        RECT 131.800 84.800 133.800 85.100 ;
        RECT 131.800 81.100 132.200 84.800 ;
        RECT 133.400 81.100 133.800 84.800 ;
        RECT 134.200 84.800 135.500 85.100 ;
        RECT 134.200 81.100 134.600 84.800 ;
        RECT 135.800 84.600 136.300 85.100 ;
        RECT 137.400 87.700 137.800 89.900 ;
        RECT 139.500 89.200 140.100 89.900 ;
        RECT 139.500 88.900 140.200 89.200 ;
        RECT 141.800 88.900 142.200 89.900 ;
        RECT 144.000 89.200 144.400 89.900 ;
        RECT 144.000 88.900 145.000 89.200 ;
        RECT 139.800 88.500 140.200 88.900 ;
        RECT 141.900 88.600 142.200 88.900 ;
        RECT 141.900 88.300 143.300 88.600 ;
        RECT 142.900 88.200 143.300 88.300 ;
        RECT 143.800 88.200 144.200 88.600 ;
        RECT 144.600 88.500 145.000 88.900 ;
        RECT 138.900 87.700 139.300 87.800 ;
        RECT 137.400 87.400 139.300 87.700 ;
        RECT 137.400 85.700 137.800 87.400 ;
        RECT 140.900 87.100 141.300 87.200 ;
        RECT 143.800 87.100 144.100 88.200 ;
        RECT 146.200 87.500 146.600 89.900 ;
        RECT 147.000 87.900 147.400 89.900 ;
        RECT 147.800 88.000 148.200 89.900 ;
        RECT 149.400 88.000 149.800 89.900 ;
        RECT 147.800 87.900 149.800 88.000 ;
        RECT 150.200 88.500 150.600 89.500 ;
        RECT 147.100 87.200 147.400 87.900 ;
        RECT 147.900 87.700 149.700 87.900 ;
        RECT 150.200 87.400 150.500 88.500 ;
        RECT 152.300 88.000 152.700 89.500 ;
        RECT 156.700 88.200 157.100 88.600 ;
        RECT 152.300 87.700 153.100 88.000 ;
        RECT 156.600 87.800 157.000 88.200 ;
        RECT 157.400 87.900 157.800 89.900 ;
        RECT 152.700 87.500 153.100 87.700 ;
        RECT 149.000 87.200 149.400 87.400 ;
        RECT 145.400 87.100 146.200 87.200 ;
        RECT 140.700 86.800 146.200 87.100 ;
        RECT 147.000 86.800 148.300 87.200 ;
        RECT 149.000 86.900 149.800 87.200 ;
        RECT 150.200 87.100 152.300 87.400 ;
        RECT 149.400 86.800 149.800 86.900 ;
        RECT 151.800 86.900 152.300 87.100 ;
        RECT 152.800 87.200 153.100 87.500 ;
        RECT 152.800 87.100 153.800 87.200 ;
        RECT 156.600 87.100 157.000 87.200 ;
        RECT 139.800 86.400 140.200 86.500 ;
        RECT 138.300 86.100 140.200 86.400 ;
        RECT 138.300 86.000 138.700 86.100 ;
        RECT 139.100 85.700 139.500 85.800 ;
        RECT 137.400 85.400 139.500 85.700 ;
        RECT 135.800 81.100 136.200 84.600 ;
        RECT 137.400 81.100 137.800 85.400 ;
        RECT 140.700 85.200 141.000 86.800 ;
        RECT 144.300 86.700 144.700 86.800 ;
        RECT 143.800 86.200 144.200 86.300 ;
        RECT 145.100 86.200 145.500 86.300 ;
        RECT 143.000 85.900 145.500 86.200 ;
        RECT 143.000 85.800 143.400 85.900 ;
        RECT 143.800 85.500 146.600 85.600 ;
        RECT 143.700 85.400 146.600 85.500 ;
        RECT 139.800 84.900 141.000 85.200 ;
        RECT 141.700 85.300 146.600 85.400 ;
        RECT 141.700 85.100 144.100 85.300 ;
        RECT 139.800 84.400 140.100 84.900 ;
        RECT 139.400 84.000 140.100 84.400 ;
        RECT 140.900 84.500 141.300 84.600 ;
        RECT 141.700 84.500 142.000 85.100 ;
        RECT 140.900 84.200 142.000 84.500 ;
        RECT 142.300 84.500 145.000 84.800 ;
        RECT 142.300 84.400 142.700 84.500 ;
        RECT 144.600 84.400 145.000 84.500 ;
        RECT 141.500 83.700 141.900 83.800 ;
        RECT 142.900 83.700 143.300 83.800 ;
        RECT 139.800 83.100 140.200 83.500 ;
        RECT 141.500 83.400 143.300 83.700 ;
        RECT 141.900 83.100 142.200 83.400 ;
        RECT 144.600 83.100 145.000 83.500 ;
        RECT 139.500 81.100 140.100 83.100 ;
        RECT 141.800 81.100 142.200 83.100 ;
        RECT 144.000 82.800 145.000 83.100 ;
        RECT 144.000 81.100 144.400 82.800 ;
        RECT 146.200 81.100 146.600 85.300 ;
        RECT 147.000 85.100 147.400 85.200 ;
        RECT 148.000 85.100 148.300 86.800 ;
        RECT 148.600 85.800 149.000 86.600 ;
        RECT 150.200 85.800 150.600 86.600 ;
        RECT 151.000 85.800 151.400 86.600 ;
        RECT 151.800 86.500 152.500 86.900 ;
        RECT 152.800 86.800 157.000 87.100 ;
        RECT 151.800 85.500 152.100 86.500 ;
        RECT 150.200 85.200 152.100 85.500 ;
        RECT 147.000 84.800 147.700 85.100 ;
        RECT 148.000 84.800 148.500 85.100 ;
        RECT 147.400 84.200 147.700 84.800 ;
        RECT 147.400 83.800 147.800 84.200 ;
        RECT 148.100 82.200 148.500 84.800 ;
        RECT 150.200 83.500 150.500 85.200 ;
        RECT 152.800 84.900 153.100 86.800 ;
        RECT 153.400 85.400 153.800 86.200 ;
        RECT 156.600 86.100 157.000 86.200 ;
        RECT 157.500 86.100 157.800 87.900 ;
        RECT 158.200 86.400 158.600 87.200 ;
        RECT 159.000 87.100 159.400 87.200 ;
        RECT 159.800 87.100 160.200 89.900 ;
        RECT 160.600 88.100 161.000 88.600 ;
        RECT 161.400 88.100 161.800 89.900 ;
        RECT 163.500 89.200 164.100 89.900 ;
        RECT 163.500 88.900 164.200 89.200 ;
        RECT 165.800 88.900 166.200 89.900 ;
        RECT 168.000 89.200 168.400 89.900 ;
        RECT 168.000 88.900 169.000 89.200 ;
        RECT 163.800 88.500 164.200 88.900 ;
        RECT 165.900 88.600 166.200 88.900 ;
        RECT 165.900 88.300 167.300 88.600 ;
        RECT 166.900 88.200 167.300 88.300 ;
        RECT 167.800 88.200 168.200 88.600 ;
        RECT 168.600 88.500 169.000 88.900 ;
        RECT 160.600 87.800 161.800 88.100 ;
        RECT 159.000 86.800 160.200 87.100 ;
        RECT 159.000 86.100 159.400 86.200 ;
        RECT 156.600 85.800 157.800 86.100 ;
        RECT 158.600 85.800 159.400 86.100 ;
        RECT 156.700 85.100 157.000 85.800 ;
        RECT 158.600 85.600 159.000 85.800 ;
        RECT 152.300 84.600 153.100 84.900 ;
        RECT 148.100 81.800 149.000 82.200 ;
        RECT 148.100 81.100 148.500 81.800 ;
        RECT 150.200 81.500 150.600 83.500 ;
        RECT 152.300 81.100 152.700 84.600 ;
        RECT 156.600 81.100 157.000 85.100 ;
        RECT 157.400 84.800 159.400 85.100 ;
        RECT 157.400 81.100 157.800 84.800 ;
        RECT 159.000 81.100 159.400 84.800 ;
        RECT 159.800 81.100 160.200 86.800 ;
        RECT 161.400 87.700 161.800 87.800 ;
        RECT 162.900 87.700 163.300 87.800 ;
        RECT 161.400 87.400 163.300 87.700 ;
        RECT 161.400 85.700 161.800 87.400 ;
        RECT 164.900 87.100 165.300 87.200 ;
        RECT 167.800 87.100 168.100 88.200 ;
        RECT 170.200 87.500 170.600 89.900 ;
        RECT 171.000 88.000 171.400 89.900 ;
        RECT 172.600 88.000 173.000 89.900 ;
        RECT 171.000 87.900 173.000 88.000 ;
        RECT 173.400 87.900 173.800 89.900 ;
        RECT 174.500 88.200 174.900 89.900 ;
        RECT 174.500 87.900 175.400 88.200 ;
        RECT 176.600 87.900 177.000 89.900 ;
        RECT 177.400 88.000 177.800 89.900 ;
        RECT 179.000 88.000 179.400 89.900 ;
        RECT 177.400 87.900 179.400 88.000 ;
        RECT 171.100 87.700 172.900 87.900 ;
        RECT 171.400 87.200 171.800 87.400 ;
        RECT 173.400 87.200 173.700 87.900 ;
        RECT 169.400 87.100 170.200 87.200 ;
        RECT 164.700 86.800 170.200 87.100 ;
        RECT 171.000 86.900 171.800 87.200 ;
        RECT 171.000 86.800 171.400 86.900 ;
        RECT 172.500 86.800 173.800 87.200 ;
        RECT 163.800 86.400 164.200 86.500 ;
        RECT 162.300 86.100 164.200 86.400 ;
        RECT 164.700 86.200 165.000 86.800 ;
        RECT 168.300 86.700 168.700 86.800 ;
        RECT 169.100 86.200 169.500 86.300 ;
        RECT 162.300 86.000 162.700 86.100 ;
        RECT 164.600 85.800 165.000 86.200 ;
        RECT 167.000 85.900 169.500 86.200 ;
        RECT 167.000 85.800 167.400 85.900 ;
        RECT 171.800 85.800 172.200 86.600 ;
        RECT 163.100 85.700 163.500 85.800 ;
        RECT 161.400 85.400 163.500 85.700 ;
        RECT 161.400 81.100 161.800 85.400 ;
        RECT 164.700 85.200 165.000 85.800 ;
        RECT 167.800 85.500 170.600 85.600 ;
        RECT 167.700 85.400 170.600 85.500 ;
        RECT 163.800 84.900 165.000 85.200 ;
        RECT 165.700 85.300 170.600 85.400 ;
        RECT 165.700 85.100 168.100 85.300 ;
        RECT 163.800 84.400 164.100 84.900 ;
        RECT 163.400 84.000 164.100 84.400 ;
        RECT 164.900 84.500 165.300 84.600 ;
        RECT 165.700 84.500 166.000 85.100 ;
        RECT 164.900 84.200 166.000 84.500 ;
        RECT 166.300 84.500 169.000 84.800 ;
        RECT 166.300 84.400 166.700 84.500 ;
        RECT 168.600 84.400 169.000 84.500 ;
        RECT 165.500 83.700 165.900 83.800 ;
        RECT 166.900 83.700 167.300 83.800 ;
        RECT 163.800 83.100 164.200 83.500 ;
        RECT 165.500 83.400 167.300 83.700 ;
        RECT 165.900 83.100 166.200 83.400 ;
        RECT 168.600 83.100 169.000 83.500 ;
        RECT 163.500 81.100 164.100 83.100 ;
        RECT 165.800 81.100 166.200 83.100 ;
        RECT 168.000 82.800 169.000 83.100 ;
        RECT 168.000 81.100 168.400 82.800 ;
        RECT 170.200 81.100 170.600 85.300 ;
        RECT 172.500 85.200 172.800 86.800 ;
        RECT 171.800 84.800 172.800 85.200 ;
        RECT 173.400 85.100 173.800 85.200 ;
        RECT 173.100 84.800 173.800 85.100 ;
        RECT 172.300 81.100 172.700 84.800 ;
        RECT 173.100 84.200 173.400 84.800 ;
        RECT 174.200 84.400 174.600 85.200 ;
        RECT 175.000 85.100 175.400 87.900 ;
        RECT 175.800 86.800 176.200 87.600 ;
        RECT 176.700 87.200 177.000 87.900 ;
        RECT 177.500 87.700 179.300 87.900 ;
        RECT 179.800 87.700 180.200 89.900 ;
        RECT 181.900 89.200 182.500 89.900 ;
        RECT 181.900 88.900 182.600 89.200 ;
        RECT 184.200 88.900 184.600 89.900 ;
        RECT 186.400 89.200 186.800 89.900 ;
        RECT 186.400 88.900 187.400 89.200 ;
        RECT 182.200 88.500 182.600 88.900 ;
        RECT 184.300 88.600 184.600 88.900 ;
        RECT 184.300 88.300 185.700 88.600 ;
        RECT 185.300 88.200 185.700 88.300 ;
        RECT 186.200 88.200 186.600 88.600 ;
        RECT 187.000 88.500 187.400 88.900 ;
        RECT 181.300 87.700 181.700 87.800 ;
        RECT 179.800 87.400 181.700 87.700 ;
        RECT 178.600 87.200 179.000 87.400 ;
        RECT 176.600 86.800 177.900 87.200 ;
        RECT 178.600 86.900 179.400 87.200 ;
        RECT 179.000 86.800 179.400 86.900 ;
        RECT 176.600 86.100 177.000 86.200 ;
        RECT 177.600 86.100 177.900 86.800 ;
        RECT 176.600 85.800 177.900 86.100 ;
        RECT 178.200 85.800 178.600 86.600 ;
        RECT 176.600 85.100 177.000 85.200 ;
        RECT 177.600 85.100 177.900 85.800 ;
        RECT 179.800 85.700 180.200 87.400 ;
        RECT 183.300 87.100 183.700 87.200 ;
        RECT 186.200 87.100 186.500 88.200 ;
        RECT 188.600 87.500 189.000 89.900 ;
        RECT 191.300 88.000 191.700 89.500 ;
        RECT 193.400 88.500 193.800 89.500 ;
        RECT 190.900 87.700 191.700 88.000 ;
        RECT 190.900 87.500 191.300 87.700 ;
        RECT 190.900 87.200 191.200 87.500 ;
        RECT 193.500 87.400 193.800 88.500 ;
        RECT 187.800 87.100 188.600 87.200 ;
        RECT 189.400 87.100 189.800 87.200 ;
        RECT 183.100 86.800 189.800 87.100 ;
        RECT 190.200 86.800 191.200 87.200 ;
        RECT 191.700 87.100 193.800 87.400 ;
        RECT 191.700 86.900 192.200 87.100 ;
        RECT 182.200 86.400 182.600 86.500 ;
        RECT 180.700 86.100 182.600 86.400 ;
        RECT 183.100 86.200 183.400 86.800 ;
        RECT 186.700 86.700 187.100 86.800 ;
        RECT 187.500 86.200 187.900 86.300 ;
        RECT 190.900 86.200 191.200 86.800 ;
        RECT 191.500 86.500 192.200 86.900 ;
        RECT 180.700 86.000 181.100 86.100 ;
        RECT 183.000 85.800 183.400 86.200 ;
        RECT 185.400 85.900 187.900 86.200 ;
        RECT 185.400 85.800 185.800 85.900 ;
        RECT 181.500 85.700 181.900 85.800 ;
        RECT 179.800 85.400 181.900 85.700 ;
        RECT 175.000 84.800 177.300 85.100 ;
        RECT 177.600 84.800 178.100 85.100 ;
        RECT 173.000 83.800 173.400 84.200 ;
        RECT 175.000 81.100 175.400 84.800 ;
        RECT 177.000 84.200 177.300 84.800 ;
        RECT 177.000 83.800 177.400 84.200 ;
        RECT 177.700 81.100 178.100 84.800 ;
        RECT 179.800 81.100 180.200 85.400 ;
        RECT 183.100 85.200 183.400 85.800 ;
        RECT 186.200 85.500 189.000 85.600 ;
        RECT 186.100 85.400 189.000 85.500 ;
        RECT 190.200 85.400 190.600 86.200 ;
        RECT 190.900 85.800 191.400 86.200 ;
        RECT 182.200 84.900 183.400 85.200 ;
        RECT 184.100 85.300 189.000 85.400 ;
        RECT 184.100 85.100 186.500 85.300 ;
        RECT 182.200 84.400 182.500 84.900 ;
        RECT 181.800 84.000 182.500 84.400 ;
        RECT 183.300 84.500 183.700 84.600 ;
        RECT 184.100 84.500 184.400 85.100 ;
        RECT 183.300 84.200 184.400 84.500 ;
        RECT 184.700 84.500 187.400 84.800 ;
        RECT 184.700 84.400 185.100 84.500 ;
        RECT 187.000 84.400 187.400 84.500 ;
        RECT 183.900 83.700 184.300 83.800 ;
        RECT 185.300 83.700 185.700 83.800 ;
        RECT 182.200 83.100 182.600 83.500 ;
        RECT 183.900 83.400 185.700 83.700 ;
        RECT 184.300 83.100 184.600 83.400 ;
        RECT 187.000 83.100 187.400 83.500 ;
        RECT 181.900 81.100 182.500 83.100 ;
        RECT 184.200 81.100 184.600 83.100 ;
        RECT 186.400 82.800 187.400 83.100 ;
        RECT 186.400 81.100 186.800 82.800 ;
        RECT 188.600 81.100 189.000 85.300 ;
        RECT 190.900 84.900 191.200 85.800 ;
        RECT 191.900 85.500 192.200 86.500 ;
        RECT 192.600 85.800 193.000 86.600 ;
        RECT 193.400 85.800 193.800 86.600 ;
        RECT 191.900 85.200 193.800 85.500 ;
        RECT 190.900 84.600 191.700 84.900 ;
        RECT 191.300 81.100 191.700 84.600 ;
        RECT 193.500 83.500 193.800 85.200 ;
        RECT 193.400 81.500 193.800 83.500 ;
        RECT 194.200 81.100 194.600 89.900 ;
        RECT 195.000 88.100 195.400 88.600 ;
        RECT 195.800 88.100 196.200 89.900 ;
        RECT 197.900 89.200 198.500 89.900 ;
        RECT 197.900 88.900 198.600 89.200 ;
        RECT 200.200 88.900 200.600 89.900 ;
        RECT 202.400 89.200 202.800 89.900 ;
        RECT 202.400 88.900 203.400 89.200 ;
        RECT 198.200 88.500 198.600 88.900 ;
        RECT 200.300 88.600 200.600 88.900 ;
        RECT 200.300 88.300 201.700 88.600 ;
        RECT 201.300 88.200 201.700 88.300 ;
        RECT 202.200 88.200 202.600 88.600 ;
        RECT 203.000 88.500 203.400 88.900 ;
        RECT 195.000 87.800 196.200 88.100 ;
        RECT 195.800 87.700 196.200 87.800 ;
        RECT 197.300 87.700 197.700 87.800 ;
        RECT 195.800 87.400 197.700 87.700 ;
        RECT 195.800 85.700 196.200 87.400 ;
        RECT 202.200 87.200 202.500 88.200 ;
        RECT 204.600 87.500 205.000 89.900 ;
        RECT 199.300 87.100 199.700 87.200 ;
        RECT 201.400 87.100 201.800 87.200 ;
        RECT 202.200 87.100 202.600 87.200 ;
        RECT 203.800 87.100 204.600 87.200 ;
        RECT 199.100 86.800 204.600 87.100 ;
        RECT 198.200 86.400 198.600 86.500 ;
        RECT 196.700 86.100 198.600 86.400 ;
        RECT 196.700 86.000 197.100 86.100 ;
        RECT 197.500 85.700 197.900 85.800 ;
        RECT 195.800 85.400 197.900 85.700 ;
        RECT 195.800 81.100 196.200 85.400 ;
        RECT 199.100 85.200 199.400 86.800 ;
        RECT 202.700 86.700 203.100 86.800 ;
        RECT 203.500 86.200 203.900 86.300 ;
        RECT 201.400 85.900 203.900 86.200 ;
        RECT 201.400 85.800 201.800 85.900 ;
        RECT 202.200 85.500 205.000 85.600 ;
        RECT 202.100 85.400 205.000 85.500 ;
        RECT 198.200 84.900 199.400 85.200 ;
        RECT 200.100 85.300 205.000 85.400 ;
        RECT 200.100 85.100 202.500 85.300 ;
        RECT 198.200 84.400 198.500 84.900 ;
        RECT 197.800 84.000 198.500 84.400 ;
        RECT 199.300 84.500 199.700 84.600 ;
        RECT 200.100 84.500 200.400 85.100 ;
        RECT 199.300 84.200 200.400 84.500 ;
        RECT 200.700 84.500 203.400 84.800 ;
        RECT 200.700 84.400 201.100 84.500 ;
        RECT 203.000 84.400 203.400 84.500 ;
        RECT 199.900 83.700 200.300 83.800 ;
        RECT 201.300 83.700 201.700 83.800 ;
        RECT 198.200 83.100 198.600 83.500 ;
        RECT 199.900 83.400 201.700 83.700 ;
        RECT 200.300 83.100 200.600 83.400 ;
        RECT 203.000 83.100 203.400 83.500 ;
        RECT 197.900 81.100 198.500 83.100 ;
        RECT 200.200 81.100 200.600 83.100 ;
        RECT 202.400 82.800 203.400 83.100 ;
        RECT 202.400 81.100 202.800 82.800 ;
        RECT 204.600 81.100 205.000 85.300 ;
        RECT 0.600 75.700 1.000 79.900 ;
        RECT 2.800 78.200 3.200 79.900 ;
        RECT 2.200 77.900 3.200 78.200 ;
        RECT 5.000 77.900 5.400 79.900 ;
        RECT 7.100 77.900 7.700 79.900 ;
        RECT 2.200 77.500 2.600 77.900 ;
        RECT 5.000 77.600 5.300 77.900 ;
        RECT 3.900 77.300 5.700 77.600 ;
        RECT 7.000 77.500 7.400 77.900 ;
        RECT 3.900 77.200 4.300 77.300 ;
        RECT 5.300 77.200 5.700 77.300 ;
        RECT 2.200 76.500 2.600 76.600 ;
        RECT 4.500 76.500 4.900 76.600 ;
        RECT 2.200 76.200 4.900 76.500 ;
        RECT 5.200 76.500 6.300 76.800 ;
        RECT 5.200 75.900 5.500 76.500 ;
        RECT 5.900 76.400 6.300 76.500 ;
        RECT 7.100 76.600 7.800 77.000 ;
        RECT 7.100 76.100 7.400 76.600 ;
        RECT 3.100 75.700 5.500 75.900 ;
        RECT 0.600 75.600 5.500 75.700 ;
        RECT 6.200 75.800 7.400 76.100 ;
        RECT 0.600 75.500 3.500 75.600 ;
        RECT 0.600 75.400 3.400 75.500 ;
        RECT 3.800 75.100 4.200 75.200 ;
        RECT 4.600 75.100 5.000 75.200 ;
        RECT 1.700 74.800 5.000 75.100 ;
        RECT 1.700 74.700 2.100 74.800 ;
        RECT 2.500 74.200 2.900 74.300 ;
        RECT 6.200 74.200 6.500 75.800 ;
        RECT 9.400 75.600 9.800 79.900 ;
        RECT 11.500 76.300 11.900 79.900 ;
        RECT 11.000 75.900 11.900 76.300 ;
        RECT 12.600 75.900 13.000 79.900 ;
        RECT 13.400 76.200 13.800 79.900 ;
        RECT 15.000 76.200 15.400 79.900 ;
        RECT 16.200 76.800 16.600 77.200 ;
        RECT 16.200 76.200 16.500 76.800 ;
        RECT 16.900 76.200 17.300 79.900 ;
        RECT 13.400 75.900 15.400 76.200 ;
        RECT 15.800 75.900 16.500 76.200 ;
        RECT 16.800 75.900 17.300 76.200 ;
        RECT 7.700 75.300 9.800 75.600 ;
        RECT 7.700 75.200 8.100 75.300 ;
        RECT 8.500 74.900 8.900 75.000 ;
        RECT 7.000 74.600 8.900 74.900 ;
        RECT 7.000 74.500 7.400 74.600 ;
        RECT 1.000 73.900 6.500 74.200 ;
        RECT 1.000 73.800 1.800 73.900 ;
        RECT 0.600 71.100 1.000 73.500 ;
        RECT 3.100 73.200 3.400 73.900 ;
        RECT 5.900 73.800 6.300 73.900 ;
        RECT 9.400 73.600 9.800 75.300 ;
        RECT 11.100 74.200 11.400 75.900 ;
        RECT 11.800 74.800 12.200 75.600 ;
        RECT 12.700 75.200 13.000 75.900 ;
        RECT 15.800 75.800 16.200 75.900 ;
        RECT 14.600 75.200 15.000 75.400 ;
        RECT 12.600 74.900 13.800 75.200 ;
        RECT 14.600 74.900 15.400 75.200 ;
        RECT 12.600 74.800 13.000 74.900 ;
        RECT 11.000 73.800 11.400 74.200 ;
        RECT 7.900 73.300 9.800 73.600 ;
        RECT 7.900 73.200 8.300 73.300 ;
        RECT 2.200 72.100 2.600 72.500 ;
        RECT 3.000 72.400 3.400 73.200 ;
        RECT 9.400 73.100 9.800 73.300 ;
        RECT 10.200 73.100 10.600 73.200 ;
        RECT 11.100 73.100 11.400 73.800 ;
        RECT 12.600 73.100 13.000 73.200 ;
        RECT 13.500 73.100 13.800 74.900 ;
        RECT 15.000 74.800 15.400 74.900 ;
        RECT 15.800 75.100 16.200 75.200 ;
        RECT 16.800 75.100 17.100 75.900 ;
        RECT 19.000 75.700 19.400 79.900 ;
        RECT 21.200 78.200 21.600 79.900 ;
        RECT 20.600 77.900 21.600 78.200 ;
        RECT 23.400 77.900 23.800 79.900 ;
        RECT 25.500 77.900 26.100 79.900 ;
        RECT 20.600 77.500 21.000 77.900 ;
        RECT 23.400 77.600 23.700 77.900 ;
        RECT 22.300 77.300 24.100 77.600 ;
        RECT 25.400 77.500 25.800 77.900 ;
        RECT 22.300 77.200 22.700 77.300 ;
        RECT 23.700 77.200 24.100 77.300 ;
        RECT 20.600 76.500 21.000 76.600 ;
        RECT 22.900 76.500 23.300 76.600 ;
        RECT 20.600 76.200 23.300 76.500 ;
        RECT 23.600 76.500 24.700 76.800 ;
        RECT 23.600 75.900 23.900 76.500 ;
        RECT 24.300 76.400 24.700 76.500 ;
        RECT 25.500 76.600 26.200 77.000 ;
        RECT 25.500 76.100 25.800 76.600 ;
        RECT 21.500 75.700 23.900 75.900 ;
        RECT 19.000 75.600 23.900 75.700 ;
        RECT 24.600 75.800 25.800 76.100 ;
        RECT 19.000 75.500 21.900 75.600 ;
        RECT 19.000 75.400 21.800 75.500 ;
        RECT 15.800 74.800 17.100 75.100 ;
        RECT 14.200 73.800 14.600 74.600 ;
        RECT 16.800 74.200 17.100 74.800 ;
        RECT 17.400 75.100 17.800 75.200 ;
        RECT 18.200 75.100 18.600 75.200 ;
        RECT 22.200 75.100 22.600 75.200 ;
        RECT 17.400 74.800 18.600 75.100 ;
        RECT 20.100 74.800 22.600 75.100 ;
        RECT 17.400 74.400 17.800 74.800 ;
        RECT 20.100 74.700 20.500 74.800 ;
        RECT 21.400 74.700 21.800 74.800 ;
        RECT 20.900 74.200 21.300 74.300 ;
        RECT 24.600 74.200 24.900 75.800 ;
        RECT 27.800 75.600 28.200 79.900 ;
        RECT 26.100 75.300 28.200 75.600 ;
        RECT 26.100 75.200 26.500 75.300 ;
        RECT 26.900 74.900 27.300 75.000 ;
        RECT 25.400 74.600 27.300 74.900 ;
        RECT 25.400 74.500 25.800 74.600 ;
        RECT 15.800 73.800 17.100 74.200 ;
        RECT 18.200 74.100 18.600 74.200 ;
        RECT 17.800 73.800 18.600 74.100 ;
        RECT 19.400 73.900 24.900 74.200 ;
        RECT 19.400 73.800 20.200 73.900 ;
        RECT 15.900 73.100 16.200 73.800 ;
        RECT 17.800 73.600 18.200 73.800 ;
        RECT 16.700 73.100 18.500 73.300 ;
        RECT 9.400 72.800 10.600 73.100 ;
        RECT 11.000 72.800 13.000 73.100 ;
        RECT 3.900 72.700 4.300 72.800 ;
        RECT 3.900 72.400 5.300 72.700 ;
        RECT 5.000 72.100 5.300 72.400 ;
        RECT 7.000 72.100 7.400 72.500 ;
        RECT 2.200 71.800 3.200 72.100 ;
        RECT 2.800 71.100 3.200 71.800 ;
        RECT 5.000 71.100 5.400 72.100 ;
        RECT 7.000 71.800 7.700 72.100 ;
        RECT 7.100 71.100 7.700 71.800 ;
        RECT 9.400 71.100 9.800 72.800 ;
        RECT 10.200 72.400 10.600 72.800 ;
        RECT 11.100 72.100 11.400 72.800 ;
        RECT 12.700 72.400 13.100 72.800 ;
        RECT 11.000 71.100 11.400 72.100 ;
        RECT 13.400 71.100 13.800 73.100 ;
        RECT 15.800 71.100 16.200 73.100 ;
        RECT 16.600 73.000 18.600 73.100 ;
        RECT 16.600 71.100 17.000 73.000 ;
        RECT 18.200 71.100 18.600 73.000 ;
        RECT 19.000 71.100 19.400 73.500 ;
        RECT 21.500 73.200 21.800 73.900 ;
        RECT 24.300 73.800 24.900 73.900 ;
        RECT 20.600 72.100 21.000 72.500 ;
        RECT 21.400 72.400 21.800 73.200 ;
        RECT 24.600 73.200 24.900 73.800 ;
        RECT 27.800 73.600 28.200 75.300 ;
        RECT 26.300 73.300 28.200 73.600 ;
        RECT 28.600 73.400 29.000 74.200 ;
        RECT 26.300 73.200 26.700 73.300 ;
        RECT 24.600 72.800 25.000 73.200 ;
        RECT 22.300 72.700 22.700 72.800 ;
        RECT 22.300 72.400 23.700 72.700 ;
        RECT 23.400 72.100 23.700 72.400 ;
        RECT 25.400 72.100 25.800 72.500 ;
        RECT 20.600 71.800 21.600 72.100 ;
        RECT 21.200 71.100 21.600 71.800 ;
        RECT 23.400 71.100 23.800 72.100 ;
        RECT 25.400 71.800 26.100 72.100 ;
        RECT 25.500 71.100 26.100 71.800 ;
        RECT 27.800 71.100 28.200 73.300 ;
        RECT 29.400 73.100 29.800 79.900 ;
        RECT 30.200 75.800 30.600 76.600 ;
        RECT 29.400 72.800 30.300 73.100 ;
        RECT 29.900 72.200 30.300 72.800 ;
        RECT 29.400 71.800 30.300 72.200 ;
        RECT 29.900 71.100 30.300 71.800 ;
        RECT 31.000 71.100 31.400 79.900 ;
        RECT 32.600 75.700 33.000 79.900 ;
        RECT 34.800 78.200 35.200 79.900 ;
        RECT 34.200 77.900 35.200 78.200 ;
        RECT 37.000 77.900 37.400 79.900 ;
        RECT 39.100 77.900 39.700 79.900 ;
        RECT 34.200 77.500 34.600 77.900 ;
        RECT 37.000 77.600 37.300 77.900 ;
        RECT 35.900 77.300 37.700 77.600 ;
        RECT 39.000 77.500 39.400 77.900 ;
        RECT 35.900 77.200 36.300 77.300 ;
        RECT 37.300 77.200 37.700 77.300 ;
        RECT 41.400 77.100 41.800 79.900 ;
        RECT 42.200 77.100 42.600 77.200 ;
        RECT 34.200 76.500 34.600 76.600 ;
        RECT 36.500 76.500 36.900 76.600 ;
        RECT 34.200 76.200 36.900 76.500 ;
        RECT 37.200 76.500 38.300 76.800 ;
        RECT 37.200 75.900 37.500 76.500 ;
        RECT 37.900 76.400 38.300 76.500 ;
        RECT 39.100 76.600 39.800 77.000 ;
        RECT 41.400 76.800 42.600 77.100 ;
        RECT 39.100 76.100 39.400 76.600 ;
        RECT 35.100 75.700 37.500 75.900 ;
        RECT 32.600 75.600 37.500 75.700 ;
        RECT 38.200 75.800 39.400 76.100 ;
        RECT 32.600 75.500 35.500 75.600 ;
        RECT 32.600 75.400 35.400 75.500 ;
        RECT 35.800 75.100 36.200 75.200 ;
        RECT 33.700 74.800 36.200 75.100 ;
        RECT 33.700 74.700 34.100 74.800 ;
        RECT 34.500 74.200 34.900 74.300 ;
        RECT 38.200 74.200 38.500 75.800 ;
        RECT 41.400 75.600 41.800 76.800 ;
        RECT 39.700 75.300 41.800 75.600 ;
        RECT 39.700 75.200 40.100 75.300 ;
        RECT 40.500 74.900 40.900 75.000 ;
        RECT 39.000 74.600 40.900 74.900 ;
        RECT 39.000 74.500 39.400 74.600 ;
        RECT 33.000 73.900 38.500 74.200 ;
        RECT 33.000 73.800 33.800 73.900 ;
        RECT 31.800 72.400 32.200 73.200 ;
        RECT 32.600 71.100 33.000 73.500 ;
        RECT 35.100 72.800 35.400 73.900 ;
        RECT 36.600 73.800 37.000 73.900 ;
        RECT 37.900 73.800 38.300 73.900 ;
        RECT 41.400 73.600 41.800 75.300 ;
        RECT 43.000 75.100 43.400 79.900 ;
        RECT 45.000 76.800 45.400 77.200 ;
        RECT 43.800 75.800 44.200 76.600 ;
        RECT 45.000 76.200 45.300 76.800 ;
        RECT 45.700 76.200 46.100 79.900 ;
        RECT 44.600 75.900 45.300 76.200 ;
        RECT 45.600 75.900 46.100 76.200 ;
        RECT 49.100 76.200 49.500 79.900 ;
        RECT 53.900 78.200 54.300 79.900 ;
        RECT 53.400 77.800 54.300 78.200 ;
        RECT 49.800 76.800 50.200 77.200 ;
        RECT 49.900 76.200 50.200 76.800 ;
        RECT 53.900 76.200 54.300 77.800 ;
        RECT 54.600 76.800 55.000 77.200 ;
        RECT 54.700 76.200 55.000 76.800 ;
        RECT 56.600 76.400 57.000 79.900 ;
        RECT 49.100 75.900 49.600 76.200 ;
        RECT 49.900 76.100 50.600 76.200 ;
        RECT 49.900 75.900 51.300 76.100 ;
        RECT 53.900 75.900 54.400 76.200 ;
        RECT 54.700 75.900 55.400 76.200 ;
        RECT 44.600 75.800 45.000 75.900 ;
        RECT 44.600 75.100 44.900 75.800 ;
        RECT 43.000 74.800 44.900 75.100 ;
        RECT 39.900 73.300 41.800 73.600 ;
        RECT 42.200 73.400 42.600 74.200 ;
        RECT 39.900 73.200 40.300 73.300 ;
        RECT 34.200 72.100 34.600 72.500 ;
        RECT 35.000 72.400 35.400 72.800 ;
        RECT 35.900 72.700 36.300 72.800 ;
        RECT 35.900 72.400 37.300 72.700 ;
        RECT 37.000 72.100 37.300 72.400 ;
        RECT 39.000 72.100 39.400 72.500 ;
        RECT 34.200 71.800 35.200 72.100 ;
        RECT 34.800 71.100 35.200 71.800 ;
        RECT 37.000 71.100 37.400 72.100 ;
        RECT 39.000 71.800 39.700 72.100 ;
        RECT 39.100 71.100 39.700 71.800 ;
        RECT 41.400 71.100 41.800 73.300 ;
        RECT 43.000 73.100 43.400 74.800 ;
        RECT 45.600 74.200 45.900 75.900 ;
        RECT 49.300 75.200 49.600 75.900 ;
        RECT 50.200 75.800 51.300 75.900 ;
        RECT 46.200 74.400 46.600 75.200 ;
        RECT 48.600 74.400 49.000 75.200 ;
        RECT 49.300 74.800 49.800 75.200 ;
        RECT 52.600 75.100 53.000 75.200 ;
        RECT 53.400 75.100 53.800 75.200 ;
        RECT 52.600 74.800 53.800 75.100 ;
        RECT 49.300 74.200 49.600 74.800 ;
        RECT 53.400 74.400 53.800 74.800 ;
        RECT 54.100 74.200 54.400 75.900 ;
        RECT 55.000 75.800 55.400 75.900 ;
        RECT 56.500 75.900 57.000 76.400 ;
        RECT 58.200 76.200 58.600 79.900 ;
        RECT 57.300 75.900 58.600 76.200 ;
        RECT 59.300 76.300 59.700 79.900 ;
        RECT 59.300 75.900 60.200 76.300 ;
        RECT 62.700 75.900 63.700 79.900 ;
        RECT 66.700 76.200 67.100 79.900 ;
        RECT 67.400 76.800 67.800 77.200 ;
        RECT 67.500 76.200 67.800 76.800 ;
        RECT 69.900 76.200 70.300 79.900 ;
        RECT 73.100 79.200 74.100 79.900 ;
        RECT 72.600 78.800 74.100 79.200 ;
        RECT 70.600 76.800 71.000 77.200 ;
        RECT 70.700 76.200 71.000 76.800 ;
        RECT 66.700 75.900 67.200 76.200 ;
        RECT 67.500 75.900 68.200 76.200 ;
        RECT 69.900 75.900 70.400 76.200 ;
        RECT 70.700 75.900 71.400 76.200 ;
        RECT 73.100 75.900 74.100 78.800 ;
        RECT 77.100 75.900 78.100 79.900 ;
        RECT 81.100 75.900 82.100 79.900 ;
        RECT 85.100 76.200 85.500 79.900 ;
        RECT 85.800 76.800 86.200 77.200 ;
        RECT 85.900 76.200 86.200 76.800 ;
        RECT 85.100 75.900 85.600 76.200 ;
        RECT 85.900 75.900 86.600 76.200 ;
        RECT 87.000 75.900 87.400 79.900 ;
        RECT 87.800 76.200 88.200 79.900 ;
        RECT 89.400 76.200 89.800 79.900 ;
        RECT 87.800 75.900 89.800 76.200 ;
        RECT 91.500 75.900 92.500 79.900 ;
        RECT 95.500 76.300 95.900 79.900 ;
        RECT 95.000 75.900 95.900 76.300 ;
        RECT 55.000 75.100 55.300 75.800 ;
        RECT 55.000 74.800 56.100 75.100 ;
        RECT 43.800 74.100 44.200 74.200 ;
        RECT 44.600 74.100 45.900 74.200 ;
        RECT 47.000 74.100 47.400 74.200 ;
        RECT 43.800 73.800 45.900 74.100 ;
        RECT 46.600 73.800 47.400 74.100 ;
        RECT 47.800 74.100 48.200 74.200 ;
        RECT 47.800 73.800 48.600 74.100 ;
        RECT 49.300 73.800 50.600 74.200 ;
        RECT 51.000 74.100 51.400 74.200 ;
        RECT 52.600 74.100 53.000 74.200 ;
        RECT 51.000 73.800 53.400 74.100 ;
        RECT 54.100 73.800 55.400 74.200 ;
        RECT 55.800 74.100 56.100 74.800 ;
        RECT 56.500 74.200 56.800 75.900 ;
        RECT 57.300 74.900 57.600 75.900 ;
        RECT 57.100 74.500 57.600 74.900 ;
        RECT 56.500 74.100 57.000 74.200 ;
        RECT 55.800 73.800 57.000 74.100 ;
        RECT 44.700 73.100 45.000 73.800 ;
        RECT 46.600 73.600 47.000 73.800 ;
        RECT 48.200 73.600 48.600 73.800 ;
        RECT 45.500 73.100 47.300 73.300 ;
        RECT 47.900 73.100 49.700 73.300 ;
        RECT 50.200 73.100 50.500 73.800 ;
        RECT 53.000 73.600 53.400 73.800 ;
        RECT 52.700 73.100 54.500 73.300 ;
        RECT 55.000 73.100 55.300 73.800 ;
        RECT 56.500 73.100 56.800 73.800 ;
        RECT 57.300 73.700 57.600 74.500 ;
        RECT 58.100 74.800 58.600 75.200 ;
        RECT 59.000 74.800 59.400 75.600 ;
        RECT 59.800 75.100 60.100 75.900 ;
        RECT 59.800 74.800 60.900 75.100 ;
        RECT 58.100 74.400 58.500 74.800 ;
        RECT 59.800 74.200 60.100 74.800 ;
        RECT 60.600 74.200 60.900 74.800 ;
        RECT 59.800 73.800 60.200 74.200 ;
        RECT 60.600 73.800 61.000 74.200 ;
        RECT 61.400 73.800 61.800 74.600 ;
        RECT 62.200 74.400 62.600 75.200 ;
        RECT 63.100 74.200 63.400 75.900 ;
        RECT 63.800 75.100 64.200 75.200 ;
        RECT 65.400 75.100 65.800 75.200 ;
        RECT 63.800 74.800 65.800 75.100 ;
        RECT 63.800 74.400 64.200 74.800 ;
        RECT 66.200 74.400 66.600 75.200 ;
        RECT 66.900 74.200 67.200 75.900 ;
        RECT 67.800 75.800 68.200 75.900 ;
        RECT 67.800 75.100 68.200 75.200 ;
        RECT 69.400 75.100 69.800 75.200 ;
        RECT 67.800 74.800 69.800 75.100 ;
        RECT 69.400 74.400 69.800 74.800 ;
        RECT 70.100 74.200 70.400 75.900 ;
        RECT 71.000 75.800 71.400 75.900 ;
        RECT 71.000 74.800 71.400 75.200 ;
        RECT 71.000 74.200 71.300 74.800 ;
        RECT 63.000 74.100 63.400 74.200 ;
        RECT 64.600 74.100 65.000 74.200 ;
        RECT 62.200 73.800 63.400 74.100 ;
        RECT 64.200 73.800 65.000 74.100 ;
        RECT 65.400 74.100 65.800 74.200 ;
        RECT 65.400 73.800 66.200 74.100 ;
        RECT 66.900 73.800 68.200 74.200 ;
        RECT 68.600 74.100 69.000 74.200 ;
        RECT 68.600 73.800 69.400 74.100 ;
        RECT 70.100 73.800 71.400 74.200 ;
        RECT 71.800 73.800 72.200 74.600 ;
        RECT 72.600 74.400 73.000 75.200 ;
        RECT 73.500 74.200 73.800 75.900 ;
        RECT 74.200 74.400 74.600 75.200 ;
        RECT 73.400 74.100 73.800 74.200 ;
        RECT 75.000 74.100 75.400 74.200 ;
        RECT 72.600 73.800 73.800 74.100 ;
        RECT 74.600 73.800 75.400 74.100 ;
        RECT 75.800 73.800 76.200 74.600 ;
        RECT 76.600 74.400 77.000 75.200 ;
        RECT 77.500 74.200 77.800 75.900 ;
        RECT 78.200 74.400 78.600 75.200 ;
        RECT 77.400 74.100 77.800 74.200 ;
        RECT 79.000 74.100 79.400 74.200 ;
        RECT 76.600 73.800 77.800 74.100 ;
        RECT 78.600 73.800 79.400 74.100 ;
        RECT 79.800 73.800 80.200 74.600 ;
        RECT 80.600 74.400 81.000 75.200 ;
        RECT 81.500 74.200 81.800 75.900 ;
        RECT 82.200 74.400 82.600 75.200 ;
        RECT 83.800 75.100 84.200 75.200 ;
        RECT 84.600 75.100 85.000 75.200 ;
        RECT 83.800 74.800 85.000 75.100 ;
        RECT 84.600 74.400 85.000 74.800 ;
        RECT 85.300 74.200 85.600 75.900 ;
        RECT 86.200 75.800 86.600 75.900 ;
        RECT 87.100 75.200 87.400 75.900 ;
        RECT 89.000 75.200 89.400 75.400 ;
        RECT 87.000 74.900 88.200 75.200 ;
        RECT 89.000 74.900 89.800 75.200 ;
        RECT 87.000 74.800 87.400 74.900 ;
        RECT 81.400 74.100 81.800 74.200 ;
        RECT 83.000 74.100 83.400 74.200 ;
        RECT 80.600 73.800 81.800 74.100 ;
        RECT 82.600 73.800 83.400 74.100 ;
        RECT 83.800 74.100 84.200 74.200 ;
        RECT 83.800 73.800 84.600 74.100 ;
        RECT 85.300 73.800 86.600 74.200 ;
        RECT 57.300 73.400 58.600 73.700 ;
        RECT 43.000 72.800 43.900 73.100 ;
        RECT 43.500 71.100 43.900 72.800 ;
        RECT 44.600 71.100 45.000 73.100 ;
        RECT 45.400 73.000 47.400 73.100 ;
        RECT 45.400 71.100 45.800 73.000 ;
        RECT 47.000 71.100 47.400 73.000 ;
        RECT 47.800 73.000 49.800 73.100 ;
        RECT 47.800 71.100 48.200 73.000 ;
        RECT 49.400 71.100 49.800 73.000 ;
        RECT 50.200 71.100 50.600 73.100 ;
        RECT 52.600 73.000 54.600 73.100 ;
        RECT 52.600 71.100 53.000 73.000 ;
        RECT 54.200 71.100 54.600 73.000 ;
        RECT 55.000 71.100 55.400 73.100 ;
        RECT 56.500 72.800 57.000 73.100 ;
        RECT 56.600 71.100 57.000 72.800 ;
        RECT 58.200 71.100 58.600 73.400 ;
        RECT 59.800 72.100 60.100 73.800 ;
        RECT 60.600 72.400 61.000 73.200 ;
        RECT 62.200 73.100 62.500 73.800 ;
        RECT 64.200 73.600 64.600 73.800 ;
        RECT 65.800 73.600 66.200 73.800 ;
        RECT 63.100 73.100 64.900 73.300 ;
        RECT 65.500 73.100 67.300 73.300 ;
        RECT 67.800 73.200 68.100 73.800 ;
        RECT 69.000 73.600 69.400 73.800 ;
        RECT 59.800 71.100 60.200 72.100 ;
        RECT 61.400 71.400 61.800 73.100 ;
        RECT 62.200 71.700 62.600 73.100 ;
        RECT 63.000 73.000 65.000 73.100 ;
        RECT 63.000 71.400 63.400 73.000 ;
        RECT 61.400 71.100 63.400 71.400 ;
        RECT 64.600 71.100 65.000 73.000 ;
        RECT 65.400 73.000 67.400 73.100 ;
        RECT 65.400 71.100 65.800 73.000 ;
        RECT 67.000 71.100 67.400 73.000 ;
        RECT 67.800 71.100 68.200 73.200 ;
        RECT 68.700 73.100 70.500 73.300 ;
        RECT 71.000 73.100 71.300 73.800 ;
        RECT 72.600 73.100 72.900 73.800 ;
        RECT 74.600 73.600 75.000 73.800 ;
        RECT 73.500 73.100 75.300 73.300 ;
        RECT 76.600 73.100 76.900 73.800 ;
        RECT 78.600 73.600 79.000 73.800 ;
        RECT 77.500 73.100 79.300 73.300 ;
        RECT 80.600 73.100 80.900 73.800 ;
        RECT 82.600 73.600 83.000 73.800 ;
        RECT 84.200 73.600 84.600 73.800 ;
        RECT 81.500 73.100 83.300 73.300 ;
        RECT 83.900 73.100 85.700 73.300 ;
        RECT 86.200 73.100 86.500 73.800 ;
        RECT 87.000 73.100 87.400 73.200 ;
        RECT 87.900 73.100 88.200 74.900 ;
        RECT 89.400 74.800 89.800 74.900 ;
        RECT 88.600 73.800 89.000 74.600 ;
        RECT 91.000 74.400 91.400 75.200 ;
        RECT 91.800 74.200 92.100 75.900 ;
        RECT 92.600 74.400 93.000 75.200 ;
        RECT 90.200 74.100 90.600 74.200 ;
        RECT 91.800 74.100 92.200 74.200 ;
        RECT 90.200 73.800 91.000 74.100 ;
        RECT 91.800 73.800 93.000 74.100 ;
        RECT 93.400 73.800 93.800 74.600 ;
        RECT 95.100 74.200 95.400 75.900 ;
        RECT 96.600 75.600 97.000 79.900 ;
        RECT 98.700 77.900 99.300 79.900 ;
        RECT 101.000 77.900 101.400 79.900 ;
        RECT 103.200 78.200 103.600 79.900 ;
        RECT 103.200 77.900 104.200 78.200 ;
        RECT 99.000 77.500 99.400 77.900 ;
        RECT 101.100 77.600 101.400 77.900 ;
        RECT 100.700 77.300 102.500 77.600 ;
        RECT 103.800 77.500 104.200 77.900 ;
        RECT 100.700 77.200 101.100 77.300 ;
        RECT 102.100 77.200 102.500 77.300 ;
        RECT 98.600 76.600 99.300 77.000 ;
        RECT 99.000 76.100 99.300 76.600 ;
        RECT 100.100 76.500 101.200 76.800 ;
        RECT 100.100 76.400 100.500 76.500 ;
        RECT 99.000 75.800 100.200 76.100 ;
        RECT 95.800 74.800 96.200 75.600 ;
        RECT 96.600 75.300 98.700 75.600 ;
        RECT 95.000 73.800 95.400 74.200 ;
        RECT 90.600 73.600 91.000 73.800 ;
        RECT 90.300 73.100 92.100 73.300 ;
        RECT 92.700 73.100 93.000 73.800 ;
        RECT 68.600 73.000 70.600 73.100 ;
        RECT 68.600 71.100 69.000 73.000 ;
        RECT 70.200 71.100 70.600 73.000 ;
        RECT 71.000 71.100 71.400 73.100 ;
        RECT 71.800 71.400 72.200 73.100 ;
        RECT 72.600 71.700 73.000 73.100 ;
        RECT 73.400 73.000 75.400 73.100 ;
        RECT 73.400 71.400 73.800 73.000 ;
        RECT 71.800 71.100 73.800 71.400 ;
        RECT 75.000 71.100 75.400 73.000 ;
        RECT 75.800 71.400 76.200 73.100 ;
        RECT 76.600 71.700 77.000 73.100 ;
        RECT 77.400 73.000 79.400 73.100 ;
        RECT 77.400 71.400 77.800 73.000 ;
        RECT 75.800 71.100 77.800 71.400 ;
        RECT 79.000 71.100 79.400 73.000 ;
        RECT 79.800 71.400 80.200 73.100 ;
        RECT 80.600 71.700 81.000 73.100 ;
        RECT 81.400 73.000 83.400 73.100 ;
        RECT 81.400 71.400 81.800 73.000 ;
        RECT 79.800 71.100 81.800 71.400 ;
        RECT 83.000 71.100 83.400 73.000 ;
        RECT 83.800 73.000 85.800 73.100 ;
        RECT 83.800 71.100 84.200 73.000 ;
        RECT 85.400 71.100 85.800 73.000 ;
        RECT 86.200 72.800 87.400 73.100 ;
        RECT 86.200 71.100 86.600 72.800 ;
        RECT 87.100 72.400 87.500 72.800 ;
        RECT 87.800 71.100 88.200 73.100 ;
        RECT 90.200 73.000 92.200 73.100 ;
        RECT 90.200 71.100 90.600 73.000 ;
        RECT 91.800 71.400 92.200 73.000 ;
        RECT 92.600 71.700 93.000 73.100 ;
        RECT 93.400 71.400 93.800 73.100 ;
        RECT 94.200 72.400 94.600 73.200 ;
        RECT 95.100 73.100 95.400 73.800 ;
        RECT 96.600 73.600 97.000 75.300 ;
        RECT 98.300 75.200 98.700 75.300 ;
        RECT 97.500 74.900 97.900 75.000 ;
        RECT 97.500 74.600 99.400 74.900 ;
        RECT 99.000 74.500 99.400 74.600 ;
        RECT 99.900 74.200 100.200 75.800 ;
        RECT 100.900 75.900 101.200 76.500 ;
        RECT 101.500 76.500 101.900 76.600 ;
        RECT 103.800 76.500 104.200 76.600 ;
        RECT 101.500 76.200 104.200 76.500 ;
        RECT 100.900 75.700 103.300 75.900 ;
        RECT 105.400 75.700 105.800 79.900 ;
        RECT 100.900 75.600 105.800 75.700 ;
        RECT 102.900 75.500 105.800 75.600 ;
        RECT 103.000 75.400 105.800 75.500 ;
        RECT 102.200 75.100 102.600 75.200 ;
        RECT 108.600 75.100 109.000 79.900 ;
        RECT 110.600 76.800 111.000 77.200 ;
        RECT 109.400 75.800 109.800 76.600 ;
        RECT 110.600 76.200 110.900 76.800 ;
        RECT 111.300 76.200 111.700 79.900 ;
        RECT 114.700 79.200 115.100 79.900 ;
        RECT 114.200 78.800 115.100 79.200 ;
        RECT 114.700 76.300 115.100 78.800 ;
        RECT 110.200 75.900 110.900 76.200 ;
        RECT 111.200 75.900 111.700 76.200 ;
        RECT 114.200 75.900 115.100 76.300 ;
        RECT 116.200 76.800 116.600 77.200 ;
        RECT 116.200 76.200 116.500 76.800 ;
        RECT 116.900 76.200 117.300 79.900 ;
        RECT 115.800 75.900 116.500 76.200 ;
        RECT 116.800 75.900 117.300 76.200 ;
        RECT 110.200 75.800 110.600 75.900 ;
        RECT 110.200 75.100 110.500 75.800 ;
        RECT 102.200 74.800 104.700 75.100 ;
        RECT 104.300 74.700 104.700 74.800 ;
        RECT 108.600 74.800 110.500 75.100 ;
        RECT 103.500 74.200 103.900 74.300 ;
        RECT 98.200 73.600 98.600 74.200 ;
        RECT 99.800 73.900 105.400 74.200 ;
        RECT 99.800 73.800 100.500 73.900 ;
        RECT 96.600 73.300 98.600 73.600 ;
        RECT 95.800 73.100 96.200 73.200 ;
        RECT 95.000 72.800 96.200 73.100 ;
        RECT 95.100 72.100 95.400 72.800 ;
        RECT 91.800 71.100 93.800 71.400 ;
        RECT 95.000 71.100 95.400 72.100 ;
        RECT 96.600 71.100 97.000 73.300 ;
        RECT 98.100 73.200 98.500 73.300 ;
        RECT 103.000 72.800 103.300 73.900 ;
        RECT 104.600 73.800 105.400 73.900 ;
        RECT 102.100 72.700 102.500 72.800 ;
        RECT 99.000 72.100 99.400 72.500 ;
        RECT 101.100 72.400 102.500 72.700 ;
        RECT 103.000 72.400 103.400 72.800 ;
        RECT 101.100 72.100 101.400 72.400 ;
        RECT 103.800 72.100 104.200 72.500 ;
        RECT 98.700 71.800 99.400 72.100 ;
        RECT 98.700 71.100 99.300 71.800 ;
        RECT 101.000 71.100 101.400 72.100 ;
        RECT 103.200 71.800 104.200 72.100 ;
        RECT 103.200 71.100 103.600 71.800 ;
        RECT 105.400 71.100 105.800 73.500 ;
        RECT 107.800 73.400 108.200 74.200 ;
        RECT 108.600 73.100 109.000 74.800 ;
        RECT 111.200 74.200 111.500 75.900 ;
        RECT 111.800 74.400 112.200 75.200 ;
        RECT 114.300 74.200 114.600 75.900 ;
        RECT 115.800 75.800 116.200 75.900 ;
        RECT 115.000 74.800 115.400 75.600 ;
        RECT 115.800 75.100 116.200 75.200 ;
        RECT 116.800 75.100 117.100 75.900 ;
        RECT 119.000 75.600 119.400 79.900 ;
        RECT 121.100 77.900 121.700 79.900 ;
        RECT 123.400 77.900 123.800 79.900 ;
        RECT 125.600 78.200 126.000 79.900 ;
        RECT 125.600 77.900 126.600 78.200 ;
        RECT 121.400 77.500 121.800 77.900 ;
        RECT 123.500 77.600 123.800 77.900 ;
        RECT 123.100 77.300 124.900 77.600 ;
        RECT 126.200 77.500 126.600 77.900 ;
        RECT 123.100 77.200 123.500 77.300 ;
        RECT 124.500 77.200 124.900 77.300 ;
        RECT 121.000 76.600 121.700 77.000 ;
        RECT 121.400 76.100 121.700 76.600 ;
        RECT 122.500 76.500 123.600 76.800 ;
        RECT 122.500 76.400 122.900 76.500 ;
        RECT 121.400 75.800 122.600 76.100 ;
        RECT 119.000 75.300 121.100 75.600 ;
        RECT 115.800 74.800 117.100 75.100 ;
        RECT 116.800 74.200 117.100 74.800 ;
        RECT 117.400 75.100 117.800 75.200 ;
        RECT 119.000 75.100 119.400 75.300 ;
        RECT 120.700 75.200 121.100 75.300 ;
        RECT 122.300 75.200 122.600 75.800 ;
        RECT 123.300 75.900 123.600 76.500 ;
        RECT 123.900 76.500 124.300 76.600 ;
        RECT 126.200 76.500 126.600 76.600 ;
        RECT 123.900 76.200 126.600 76.500 ;
        RECT 123.300 75.700 125.700 75.900 ;
        RECT 127.800 75.700 128.200 79.900 ;
        RECT 129.900 76.300 130.300 79.900 ;
        RECT 132.300 76.300 132.700 79.900 ;
        RECT 129.400 75.900 130.300 76.300 ;
        RECT 131.800 75.900 132.700 76.300 ;
        RECT 133.400 75.900 133.800 79.900 ;
        RECT 134.200 76.200 134.600 79.900 ;
        RECT 135.800 76.200 136.200 79.900 ;
        RECT 134.200 75.900 136.200 76.200 ;
        RECT 137.900 76.200 138.300 79.900 ;
        RECT 138.600 76.800 139.000 77.200 ;
        RECT 138.700 76.200 139.000 76.800 ;
        RECT 137.900 75.900 138.400 76.200 ;
        RECT 138.700 75.900 139.400 76.200 ;
        RECT 123.300 75.600 128.200 75.700 ;
        RECT 125.300 75.500 128.200 75.600 ;
        RECT 125.400 75.400 128.200 75.500 ;
        RECT 117.400 74.800 119.400 75.100 ;
        RECT 117.400 74.400 117.800 74.800 ;
        RECT 110.200 73.800 111.500 74.200 ;
        RECT 112.600 74.100 113.000 74.200 ;
        RECT 112.200 73.800 113.000 74.100 ;
        RECT 114.200 73.800 114.600 74.200 ;
        RECT 115.800 73.800 117.100 74.200 ;
        RECT 118.200 74.100 118.600 74.200 ;
        RECT 117.800 73.800 118.600 74.100 ;
        RECT 110.300 73.200 110.600 73.800 ;
        RECT 112.200 73.600 112.600 73.800 ;
        RECT 108.600 72.800 109.500 73.100 ;
        RECT 109.100 71.100 109.500 72.800 ;
        RECT 110.200 71.100 110.600 73.200 ;
        RECT 111.100 73.100 112.900 73.300 ;
        RECT 111.000 73.000 113.000 73.100 ;
        RECT 111.000 71.100 111.400 73.000 ;
        RECT 112.600 71.100 113.000 73.000 ;
        RECT 113.400 72.400 113.800 73.200 ;
        RECT 114.300 72.100 114.600 73.800 ;
        RECT 115.900 73.100 116.200 73.800 ;
        RECT 117.800 73.600 118.200 73.800 ;
        RECT 119.000 73.600 119.400 74.800 ;
        RECT 119.900 74.900 120.300 75.000 ;
        RECT 119.900 74.600 121.800 74.900 ;
        RECT 122.200 74.800 122.600 75.200 ;
        RECT 124.600 75.100 125.000 75.200 ;
        RECT 124.600 74.800 127.100 75.100 ;
        RECT 121.400 74.500 121.800 74.600 ;
        RECT 122.300 74.200 122.600 74.800 ;
        RECT 125.400 74.700 125.800 74.800 ;
        RECT 126.700 74.700 127.100 74.800 ;
        RECT 125.900 74.200 126.300 74.300 ;
        RECT 129.500 74.200 129.800 75.900 ;
        RECT 130.200 74.800 130.600 75.600 ;
        RECT 131.900 74.200 132.200 75.900 ;
        RECT 132.600 74.800 133.000 75.600 ;
        RECT 133.500 75.200 133.800 75.900 ;
        RECT 135.400 75.200 135.800 75.400 ;
        RECT 133.400 74.900 134.600 75.200 ;
        RECT 135.400 74.900 136.200 75.200 ;
        RECT 133.400 74.800 133.800 74.900 ;
        RECT 122.300 73.900 127.800 74.200 ;
        RECT 122.500 73.800 122.900 73.900 ;
        RECT 124.600 73.800 125.000 73.900 ;
        RECT 119.000 73.300 120.900 73.600 ;
        RECT 116.700 73.100 118.500 73.300 ;
        RECT 114.200 71.100 114.600 72.100 ;
        RECT 115.800 71.100 116.200 73.100 ;
        RECT 116.600 73.000 118.600 73.100 ;
        RECT 116.600 71.100 117.000 73.000 ;
        RECT 118.200 71.100 118.600 73.000 ;
        RECT 119.000 71.100 119.400 73.300 ;
        RECT 120.500 73.200 120.900 73.300 ;
        RECT 125.400 72.800 125.700 73.900 ;
        RECT 127.000 73.800 127.800 73.900 ;
        RECT 128.600 73.800 129.000 74.200 ;
        RECT 129.400 73.800 129.800 74.200 ;
        RECT 131.800 73.800 132.200 74.200 ;
        RECT 124.500 72.700 124.900 72.800 ;
        RECT 121.400 72.100 121.800 72.500 ;
        RECT 123.500 72.400 124.900 72.700 ;
        RECT 125.400 72.400 125.800 72.800 ;
        RECT 123.500 72.100 123.800 72.400 ;
        RECT 126.200 72.100 126.600 72.500 ;
        RECT 121.100 71.800 121.800 72.100 ;
        RECT 121.100 71.100 121.700 71.800 ;
        RECT 123.400 71.100 123.800 72.100 ;
        RECT 125.600 71.800 126.600 72.100 ;
        RECT 125.600 71.100 126.000 71.800 ;
        RECT 127.800 71.100 128.200 73.500 ;
        RECT 128.600 73.200 128.900 73.800 ;
        RECT 128.600 72.400 129.000 73.200 ;
        RECT 129.500 72.200 129.800 73.800 ;
        RECT 131.000 72.400 131.400 73.200 ;
        RECT 131.900 73.100 132.200 73.800 ;
        RECT 134.300 73.200 134.600 74.900 ;
        RECT 135.800 74.800 136.200 74.900 ;
        RECT 135.000 73.800 135.400 74.600 ;
        RECT 137.400 74.400 137.800 75.200 ;
        RECT 138.100 74.200 138.400 75.900 ;
        RECT 139.000 75.800 139.400 75.900 ;
        RECT 139.800 75.800 140.200 76.600 ;
        RECT 139.000 75.100 139.300 75.800 ;
        RECT 140.600 75.100 141.000 79.900 ;
        RECT 142.200 75.700 142.600 79.900 ;
        RECT 144.400 78.200 144.800 79.900 ;
        RECT 143.800 77.900 144.800 78.200 ;
        RECT 146.600 77.900 147.000 79.900 ;
        RECT 148.700 77.900 149.300 79.900 ;
        RECT 143.800 77.500 144.200 77.900 ;
        RECT 146.600 77.600 146.900 77.900 ;
        RECT 145.500 77.300 147.300 77.600 ;
        RECT 148.600 77.500 149.000 77.900 ;
        RECT 145.500 77.200 145.900 77.300 ;
        RECT 146.900 77.200 147.300 77.300 ;
        RECT 143.800 76.500 144.200 76.600 ;
        RECT 146.100 76.500 146.500 76.600 ;
        RECT 143.800 76.200 146.500 76.500 ;
        RECT 146.800 76.500 147.900 76.800 ;
        RECT 146.800 75.900 147.100 76.500 ;
        RECT 147.500 76.400 147.900 76.500 ;
        RECT 148.700 76.600 149.400 77.000 ;
        RECT 148.700 76.100 149.000 76.600 ;
        RECT 144.700 75.700 147.100 75.900 ;
        RECT 142.200 75.600 147.100 75.700 ;
        RECT 147.800 75.800 149.000 76.100 ;
        RECT 142.200 75.500 145.100 75.600 ;
        RECT 142.200 75.400 145.000 75.500 ;
        RECT 145.400 75.100 145.800 75.200 ;
        RECT 139.000 74.800 141.000 75.100 ;
        RECT 136.600 74.100 137.000 74.200 ;
        RECT 136.600 73.800 137.400 74.100 ;
        RECT 138.100 73.800 139.400 74.200 ;
        RECT 137.000 73.600 137.400 73.800 ;
        RECT 133.400 73.100 133.800 73.200 ;
        RECT 131.800 72.800 133.800 73.100 ;
        RECT 129.400 71.100 129.800 72.200 ;
        RECT 131.900 72.100 132.200 72.800 ;
        RECT 133.500 72.400 133.900 72.800 ;
        RECT 131.800 71.100 132.200 72.100 ;
        RECT 134.200 71.100 134.600 73.200 ;
        RECT 136.700 73.100 138.500 73.300 ;
        RECT 139.000 73.200 139.300 73.800 ;
        RECT 136.600 73.000 138.600 73.100 ;
        RECT 136.600 71.100 137.000 73.000 ;
        RECT 138.200 71.100 138.600 73.000 ;
        RECT 139.000 71.100 139.400 73.200 ;
        RECT 140.600 73.100 141.000 74.800 ;
        RECT 143.300 74.800 145.800 75.100 ;
        RECT 143.300 74.700 143.700 74.800 ;
        RECT 144.600 74.700 145.000 74.800 ;
        RECT 144.100 74.200 144.500 74.300 ;
        RECT 147.800 74.200 148.100 75.800 ;
        RECT 151.000 75.600 151.400 79.900 ;
        RECT 153.400 76.200 153.800 79.900 ;
        RECT 155.000 76.200 155.400 79.900 ;
        RECT 153.400 75.900 155.400 76.200 ;
        RECT 155.800 75.900 156.200 79.900 ;
        RECT 149.300 75.300 151.400 75.600 ;
        RECT 149.300 75.200 149.700 75.300 ;
        RECT 150.100 74.900 150.500 75.000 ;
        RECT 148.600 74.600 150.500 74.900 ;
        RECT 148.600 74.500 149.000 74.600 ;
        RECT 141.400 73.400 141.800 74.200 ;
        RECT 142.600 73.900 148.100 74.200 ;
        RECT 142.600 73.800 143.400 73.900 ;
        RECT 140.100 72.800 141.000 73.100 ;
        RECT 140.100 71.100 140.500 72.800 ;
        RECT 142.200 71.100 142.600 73.500 ;
        RECT 144.700 72.800 145.000 73.900 ;
        RECT 147.500 73.800 147.900 73.900 ;
        RECT 151.000 73.600 151.400 75.300 ;
        RECT 153.800 75.200 154.200 75.400 ;
        RECT 155.800 75.200 156.100 75.900 ;
        RECT 153.400 74.900 154.200 75.200 ;
        RECT 155.000 74.900 156.200 75.200 ;
        RECT 153.400 74.800 153.800 74.900 ;
        RECT 154.200 73.800 154.600 74.600 ;
        RECT 149.500 73.300 151.400 73.600 ;
        RECT 149.500 73.200 149.900 73.300 ;
        RECT 143.800 72.100 144.200 72.500 ;
        RECT 144.600 72.400 145.000 72.800 ;
        RECT 145.500 72.700 145.900 72.800 ;
        RECT 145.500 72.400 146.900 72.700 ;
        RECT 146.600 72.100 146.900 72.400 ;
        RECT 148.600 72.100 149.000 72.500 ;
        RECT 143.800 71.800 144.800 72.100 ;
        RECT 144.400 71.100 144.800 71.800 ;
        RECT 146.600 71.100 147.000 72.100 ;
        RECT 148.600 71.800 149.300 72.100 ;
        RECT 148.700 71.100 149.300 71.800 ;
        RECT 151.000 71.100 151.400 73.300 ;
        RECT 155.000 73.200 155.300 74.900 ;
        RECT 155.800 74.800 156.200 74.900 ;
        RECT 155.000 71.100 155.400 73.200 ;
        RECT 155.800 72.800 156.200 73.200 ;
        RECT 155.700 72.400 156.100 72.800 ;
        RECT 156.600 72.400 157.000 73.200 ;
        RECT 157.400 71.100 157.800 79.900 ;
        RECT 158.600 76.800 159.000 77.200 ;
        RECT 158.600 76.200 158.900 76.800 ;
        RECT 159.300 76.200 159.700 79.900 ;
        RECT 158.200 75.900 158.900 76.200 ;
        RECT 159.200 75.900 159.700 76.200 ;
        RECT 158.200 75.800 158.600 75.900 ;
        RECT 159.200 75.200 159.500 75.900 ;
        RECT 161.400 75.800 161.800 76.600 ;
        RECT 159.000 74.800 159.500 75.200 ;
        RECT 159.200 74.200 159.500 74.800 ;
        RECT 159.800 74.400 160.200 75.200 ;
        RECT 158.200 73.800 159.500 74.200 ;
        RECT 160.600 74.100 161.000 74.200 ;
        RECT 160.200 73.800 161.000 74.100 ;
        RECT 158.300 73.100 158.600 73.800 ;
        RECT 160.200 73.600 160.600 73.800 ;
        RECT 159.100 73.100 160.900 73.300 ;
        RECT 162.200 73.100 162.600 79.900 ;
        RECT 165.100 76.300 165.500 79.900 ;
        RECT 164.600 75.900 165.500 76.300 ;
        RECT 166.200 75.900 166.600 79.900 ;
        RECT 167.000 76.200 167.400 79.900 ;
        RECT 168.600 76.200 169.000 79.900 ;
        RECT 167.000 75.900 169.000 76.200 ;
        RECT 169.400 76.200 169.800 79.900 ;
        RECT 171.000 76.400 171.400 79.900 ;
        RECT 169.400 75.900 170.700 76.200 ;
        RECT 171.000 75.900 171.500 76.400 ;
        RECT 172.600 75.900 173.000 79.900 ;
        RECT 173.400 76.200 173.800 79.900 ;
        RECT 175.000 76.200 175.400 79.900 ;
        RECT 177.100 76.300 177.500 79.900 ;
        RECT 173.400 75.900 175.400 76.200 ;
        RECT 176.600 75.900 177.500 76.300 ;
        RECT 178.200 75.900 178.600 79.900 ;
        RECT 179.000 76.200 179.400 79.900 ;
        RECT 180.600 76.200 181.000 79.900 ;
        RECT 179.000 75.900 181.000 76.200 ;
        RECT 164.700 74.200 165.000 75.900 ;
        RECT 165.400 74.800 165.800 75.600 ;
        RECT 166.300 75.200 166.600 75.900 ;
        RECT 168.200 75.200 168.600 75.400 ;
        RECT 166.200 74.900 167.400 75.200 ;
        RECT 168.200 74.900 169.000 75.200 ;
        RECT 166.200 74.800 166.600 74.900 ;
        RECT 163.000 73.400 163.400 74.200 ;
        RECT 164.600 73.800 165.000 74.200 ;
        RECT 158.200 71.100 158.600 73.100 ;
        RECT 159.000 73.000 161.000 73.100 ;
        RECT 159.000 71.100 159.400 73.000 ;
        RECT 160.600 71.100 161.000 73.000 ;
        RECT 161.700 72.800 162.600 73.100 ;
        RECT 161.700 72.200 162.100 72.800 ;
        RECT 163.800 72.400 164.200 73.200 ;
        RECT 164.700 73.100 165.000 73.800 ;
        RECT 166.200 73.100 166.600 73.200 ;
        RECT 167.100 73.100 167.400 74.900 ;
        RECT 168.600 74.800 169.000 74.900 ;
        RECT 169.400 74.800 169.900 75.200 ;
        RECT 167.800 73.800 168.200 74.600 ;
        RECT 169.500 74.400 169.900 74.800 ;
        RECT 170.400 74.900 170.700 75.900 ;
        RECT 170.400 74.500 170.900 74.900 ;
        RECT 170.400 73.700 170.700 74.500 ;
        RECT 171.200 74.200 171.500 75.900 ;
        RECT 172.700 75.200 173.000 75.900 ;
        RECT 174.600 75.200 175.000 75.400 ;
        RECT 172.600 74.900 173.800 75.200 ;
        RECT 174.600 75.100 175.400 75.200 ;
        RECT 175.800 75.100 176.200 75.200 ;
        RECT 174.600 74.900 176.200 75.100 ;
        RECT 172.600 74.800 173.000 74.900 ;
        RECT 173.400 74.800 173.800 74.900 ;
        RECT 175.000 74.800 176.200 74.900 ;
        RECT 171.000 73.800 171.500 74.200 ;
        RECT 164.600 72.800 166.600 73.100 ;
        RECT 161.400 71.800 162.100 72.200 ;
        RECT 164.700 72.100 165.000 72.800 ;
        RECT 166.300 72.400 166.700 72.800 ;
        RECT 161.700 71.100 162.100 71.800 ;
        RECT 164.600 71.100 165.000 72.100 ;
        RECT 167.000 71.100 167.400 73.100 ;
        RECT 169.400 73.400 170.700 73.700 ;
        RECT 169.400 71.100 169.800 73.400 ;
        RECT 171.200 73.100 171.500 73.800 ;
        RECT 171.000 72.800 171.500 73.100 ;
        RECT 172.600 72.800 173.000 73.200 ;
        RECT 173.500 73.100 173.800 74.800 ;
        RECT 174.200 73.800 174.600 74.600 ;
        RECT 176.700 74.200 177.000 75.900 ;
        RECT 177.400 74.800 177.800 75.600 ;
        RECT 178.300 75.200 178.600 75.900 ;
        RECT 181.400 75.600 181.800 79.900 ;
        RECT 183.500 77.900 184.100 79.900 ;
        RECT 185.800 77.900 186.200 79.900 ;
        RECT 188.000 78.200 188.400 79.900 ;
        RECT 188.000 77.900 189.000 78.200 ;
        RECT 183.800 77.500 184.200 77.900 ;
        RECT 185.900 77.600 186.200 77.900 ;
        RECT 185.500 77.300 187.300 77.600 ;
        RECT 188.600 77.500 189.000 77.900 ;
        RECT 185.500 77.200 185.900 77.300 ;
        RECT 186.900 77.200 187.300 77.300 ;
        RECT 183.000 77.000 183.700 77.200 ;
        RECT 183.000 76.800 184.100 77.000 ;
        RECT 183.400 76.600 184.100 76.800 ;
        RECT 183.800 76.100 184.100 76.600 ;
        RECT 184.900 76.500 186.000 76.800 ;
        RECT 184.900 76.400 185.300 76.500 ;
        RECT 183.800 75.800 185.000 76.100 ;
        RECT 180.200 75.200 180.600 75.400 ;
        RECT 181.400 75.300 183.500 75.600 ;
        RECT 178.200 74.900 179.400 75.200 ;
        RECT 180.200 74.900 181.000 75.200 ;
        RECT 178.200 74.800 178.600 74.900 ;
        RECT 176.600 73.800 177.000 74.200 ;
        RECT 178.200 74.100 178.600 74.200 ;
        RECT 179.100 74.100 179.400 74.900 ;
        RECT 180.600 74.800 181.000 74.900 ;
        RECT 178.200 73.800 179.400 74.100 ;
        RECT 179.800 73.800 180.200 74.600 ;
        RECT 171.000 71.100 171.400 72.800 ;
        RECT 172.700 72.400 173.100 72.800 ;
        RECT 173.400 71.100 173.800 73.100 ;
        RECT 175.800 72.400 176.200 73.200 ;
        RECT 176.700 73.100 177.000 73.800 ;
        RECT 178.200 73.100 178.600 73.200 ;
        RECT 179.100 73.100 179.400 73.800 ;
        RECT 176.600 72.800 178.600 73.100 ;
        RECT 176.700 72.100 177.000 72.800 ;
        RECT 178.300 72.400 178.700 72.800 ;
        RECT 176.600 71.100 177.000 72.100 ;
        RECT 179.000 71.100 179.400 73.100 ;
        RECT 181.400 73.600 181.800 75.300 ;
        RECT 183.100 75.200 183.500 75.300 ;
        RECT 184.700 75.200 185.000 75.800 ;
        RECT 185.700 75.900 186.000 76.500 ;
        RECT 186.300 76.500 186.700 76.600 ;
        RECT 188.600 76.500 189.000 76.600 ;
        RECT 186.300 76.200 189.000 76.500 ;
        RECT 185.700 75.700 188.100 75.900 ;
        RECT 190.200 75.700 190.600 79.900 ;
        RECT 185.700 75.600 190.600 75.700 ;
        RECT 187.700 75.500 190.600 75.600 ;
        RECT 187.800 75.400 190.600 75.500 ;
        RECT 182.300 74.900 182.700 75.000 ;
        RECT 182.300 74.600 184.200 74.900 ;
        RECT 184.600 74.800 185.000 75.200 ;
        RECT 186.200 75.100 186.600 75.200 ;
        RECT 187.000 75.100 187.400 75.200 ;
        RECT 186.200 74.800 189.500 75.100 ;
        RECT 183.800 74.500 184.200 74.600 ;
        RECT 184.700 74.200 185.000 74.800 ;
        RECT 189.100 74.700 189.500 74.800 ;
        RECT 188.300 74.200 188.700 74.300 ;
        RECT 184.700 73.900 190.200 74.200 ;
        RECT 184.900 73.800 185.300 73.900 ;
        RECT 181.400 73.300 183.300 73.600 ;
        RECT 181.400 71.100 181.800 73.300 ;
        RECT 182.900 73.200 183.300 73.300 ;
        RECT 187.800 72.800 188.100 73.900 ;
        RECT 189.400 73.800 190.200 73.900 ;
        RECT 186.900 72.700 187.300 72.800 ;
        RECT 183.800 72.100 184.200 72.500 ;
        RECT 185.900 72.400 187.300 72.700 ;
        RECT 187.800 72.400 188.200 72.800 ;
        RECT 185.900 72.100 186.200 72.400 ;
        RECT 188.600 72.100 189.000 72.500 ;
        RECT 183.500 71.800 184.200 72.100 ;
        RECT 183.500 71.100 184.100 71.800 ;
        RECT 185.800 71.100 186.200 72.100 ;
        RECT 188.000 71.800 189.000 72.100 ;
        RECT 188.000 71.100 188.400 71.800 ;
        RECT 190.200 71.100 190.600 73.500 ;
        RECT 191.000 71.100 191.400 79.900 ;
        RECT 192.600 76.200 193.000 79.900 ;
        RECT 194.200 76.200 194.600 79.900 ;
        RECT 192.600 75.900 194.600 76.200 ;
        RECT 195.000 75.900 195.400 79.900 ;
        RECT 193.000 75.200 193.400 75.400 ;
        RECT 195.000 75.200 195.300 75.900 ;
        RECT 195.800 75.600 196.200 79.900 ;
        RECT 197.900 77.900 198.500 79.900 ;
        RECT 200.200 77.900 200.600 79.900 ;
        RECT 202.400 78.200 202.800 79.900 ;
        RECT 202.400 77.900 203.400 78.200 ;
        RECT 198.200 77.500 198.600 77.900 ;
        RECT 200.300 77.600 200.600 77.900 ;
        RECT 199.900 77.300 201.700 77.600 ;
        RECT 203.000 77.500 203.400 77.900 ;
        RECT 199.900 77.200 200.300 77.300 ;
        RECT 201.300 77.200 201.700 77.300 ;
        RECT 197.800 76.600 198.500 77.000 ;
        RECT 198.200 76.100 198.500 76.600 ;
        RECT 199.300 76.500 200.400 76.800 ;
        RECT 199.300 76.400 199.700 76.500 ;
        RECT 198.200 75.800 199.400 76.100 ;
        RECT 195.800 75.300 197.900 75.600 ;
        RECT 192.600 74.900 193.400 75.200 ;
        RECT 194.200 74.900 195.400 75.200 ;
        RECT 192.600 74.800 193.000 74.900 ;
        RECT 193.400 73.800 193.800 74.600 ;
        RECT 191.800 72.400 192.200 73.200 ;
        RECT 194.200 73.100 194.500 74.900 ;
        RECT 195.000 74.800 195.400 74.900 ;
        RECT 195.800 73.600 196.200 75.300 ;
        RECT 197.500 75.200 197.900 75.300 ;
        RECT 196.700 74.900 197.100 75.000 ;
        RECT 196.700 74.600 198.600 74.900 ;
        RECT 198.200 74.500 198.600 74.600 ;
        RECT 199.100 74.200 199.400 75.800 ;
        RECT 200.100 75.900 200.400 76.500 ;
        RECT 200.700 76.500 201.100 76.600 ;
        RECT 203.000 76.500 203.400 76.600 ;
        RECT 200.700 76.200 203.400 76.500 ;
        RECT 200.100 75.700 202.500 75.900 ;
        RECT 204.600 75.700 205.000 79.900 ;
        RECT 200.100 75.600 205.000 75.700 ;
        RECT 202.100 75.500 205.000 75.600 ;
        RECT 202.200 75.400 205.000 75.500 ;
        RECT 200.600 75.100 201.000 75.200 ;
        RECT 201.400 75.100 201.800 75.200 ;
        RECT 200.600 74.800 203.900 75.100 ;
        RECT 203.500 74.700 203.900 74.800 ;
        RECT 202.700 74.200 203.100 74.300 ;
        RECT 199.100 73.900 204.600 74.200 ;
        RECT 199.300 73.800 199.700 73.900 ;
        RECT 202.200 73.800 202.600 73.900 ;
        RECT 203.800 73.800 204.600 73.900 ;
        RECT 195.800 73.300 197.800 73.600 ;
        RECT 194.200 71.100 194.600 73.100 ;
        RECT 195.000 72.800 195.400 73.200 ;
        RECT 194.900 72.400 195.300 72.800 ;
        RECT 195.800 71.100 196.200 73.300 ;
        RECT 197.300 73.200 197.800 73.300 ;
        RECT 197.400 72.800 197.800 73.200 ;
        RECT 202.200 72.800 202.500 73.800 ;
        RECT 201.300 72.700 201.700 72.800 ;
        RECT 198.200 72.100 198.600 72.500 ;
        RECT 200.300 72.400 201.700 72.700 ;
        RECT 202.200 72.400 202.600 72.800 ;
        RECT 200.300 72.100 200.600 72.400 ;
        RECT 203.000 72.100 203.400 72.500 ;
        RECT 197.900 71.800 198.600 72.100 ;
        RECT 197.900 71.100 198.500 71.800 ;
        RECT 200.200 71.100 200.600 72.100 ;
        RECT 202.400 71.800 203.400 72.100 ;
        RECT 202.400 71.100 202.800 71.800 ;
        RECT 204.600 71.100 205.000 73.500 ;
        RECT 0.600 67.500 1.000 69.900 ;
        RECT 2.800 69.200 3.200 69.900 ;
        RECT 2.200 68.900 3.200 69.200 ;
        RECT 5.000 68.900 5.400 69.900 ;
        RECT 7.100 69.200 7.700 69.900 ;
        RECT 7.000 68.900 7.700 69.200 ;
        RECT 2.200 68.500 2.600 68.900 ;
        RECT 5.000 68.600 5.300 68.900 ;
        RECT 3.000 67.800 3.400 68.600 ;
        RECT 3.900 68.300 5.300 68.600 ;
        RECT 7.000 68.500 7.400 68.900 ;
        RECT 3.900 68.200 4.300 68.300 ;
        RECT 1.000 67.100 1.800 67.200 ;
        RECT 3.100 67.100 3.400 67.800 ;
        RECT 7.900 67.700 8.300 67.800 ;
        RECT 9.400 67.700 9.800 69.900 ;
        RECT 10.200 67.900 10.600 69.900 ;
        RECT 11.000 68.000 11.400 69.900 ;
        RECT 12.600 68.000 13.000 69.900 ;
        RECT 11.000 67.900 13.000 68.000 ;
        RECT 13.700 68.200 14.100 69.900 ;
        RECT 13.700 67.900 14.600 68.200 ;
        RECT 7.900 67.400 9.800 67.700 ;
        RECT 5.900 67.100 6.300 67.200 ;
        RECT 1.000 66.800 6.500 67.100 ;
        RECT 2.500 66.700 2.900 66.800 ;
        RECT 1.700 66.200 2.100 66.300 ;
        RECT 6.200 66.200 6.500 66.800 ;
        RECT 7.000 66.400 7.400 66.500 ;
        RECT 1.700 66.100 4.200 66.200 ;
        RECT 4.600 66.100 5.000 66.200 ;
        RECT 1.700 65.900 5.000 66.100 ;
        RECT 3.800 65.800 5.000 65.900 ;
        RECT 6.200 65.800 6.600 66.200 ;
        RECT 7.000 66.100 8.900 66.400 ;
        RECT 8.500 66.000 8.900 66.100 ;
        RECT 0.600 65.500 3.400 65.600 ;
        RECT 0.600 65.400 3.500 65.500 ;
        RECT 0.600 65.300 5.500 65.400 ;
        RECT 0.600 61.100 1.000 65.300 ;
        RECT 3.100 65.100 5.500 65.300 ;
        RECT 2.200 64.500 4.900 64.800 ;
        RECT 2.200 64.400 2.600 64.500 ;
        RECT 4.500 64.400 4.900 64.500 ;
        RECT 5.200 64.500 5.500 65.100 ;
        RECT 6.200 65.200 6.500 65.800 ;
        RECT 7.700 65.700 8.100 65.800 ;
        RECT 9.400 65.700 9.800 67.400 ;
        RECT 10.300 67.200 10.600 67.900 ;
        RECT 11.100 67.700 12.900 67.900 ;
        RECT 12.200 67.200 12.600 67.400 ;
        RECT 10.200 66.800 11.500 67.200 ;
        RECT 12.200 66.900 13.000 67.200 ;
        RECT 12.600 66.800 13.000 66.900 ;
        RECT 13.400 67.100 13.800 67.200 ;
        RECT 14.200 67.100 14.600 67.900 ;
        RECT 13.400 66.800 14.600 67.100 ;
        RECT 15.000 66.800 15.400 67.600 ;
        RECT 15.800 67.500 16.200 69.900 ;
        RECT 18.000 69.200 18.400 69.900 ;
        RECT 17.400 68.900 18.400 69.200 ;
        RECT 20.200 68.900 20.600 69.900 ;
        RECT 22.300 69.200 22.900 69.900 ;
        RECT 22.200 68.900 22.900 69.200 ;
        RECT 17.400 68.500 17.800 68.900 ;
        RECT 20.200 68.600 20.500 68.900 ;
        RECT 18.200 68.200 18.600 68.600 ;
        RECT 19.100 68.300 20.500 68.600 ;
        RECT 22.200 68.500 22.600 68.900 ;
        RECT 19.100 68.200 19.500 68.300 ;
        RECT 16.200 67.100 17.000 67.200 ;
        RECT 18.300 67.100 18.600 68.200 ;
        RECT 23.100 67.700 23.500 67.800 ;
        RECT 24.600 67.700 25.000 69.900 ;
        RECT 25.400 68.000 25.800 69.900 ;
        RECT 27.000 68.000 27.400 69.900 ;
        RECT 25.400 67.900 27.400 68.000 ;
        RECT 27.800 67.900 28.200 69.900 ;
        RECT 28.600 68.000 29.000 69.900 ;
        RECT 30.200 68.000 30.600 69.900 ;
        RECT 28.600 67.900 30.600 68.000 ;
        RECT 31.000 67.900 31.400 69.900 ;
        RECT 32.100 68.200 32.500 69.900 ;
        RECT 32.100 67.900 33.000 68.200 ;
        RECT 25.500 67.700 27.300 67.900 ;
        RECT 23.100 67.400 25.000 67.700 ;
        RECT 21.100 67.100 21.800 67.200 ;
        RECT 16.200 66.800 21.800 67.100 ;
        RECT 11.200 66.200 11.500 66.800 ;
        RECT 11.000 65.800 11.500 66.200 ;
        RECT 11.800 66.100 12.200 66.600 ;
        RECT 13.400 66.100 13.800 66.200 ;
        RECT 11.800 65.800 13.800 66.100 ;
        RECT 7.700 65.400 9.800 65.700 ;
        RECT 6.200 64.900 7.400 65.200 ;
        RECT 5.900 64.500 6.300 64.600 ;
        RECT 5.200 64.200 6.300 64.500 ;
        RECT 7.100 64.400 7.400 64.900 ;
        RECT 7.100 64.000 7.800 64.400 ;
        RECT 3.900 63.700 4.300 63.800 ;
        RECT 5.300 63.700 5.700 63.800 ;
        RECT 2.200 63.100 2.600 63.500 ;
        RECT 3.900 63.400 5.700 63.700 ;
        RECT 5.000 63.100 5.300 63.400 ;
        RECT 7.000 63.100 7.400 63.500 ;
        RECT 2.200 62.800 3.200 63.100 ;
        RECT 2.800 61.100 3.200 62.800 ;
        RECT 5.000 61.100 5.400 63.100 ;
        RECT 7.100 61.100 7.700 63.100 ;
        RECT 9.400 61.100 9.800 65.400 ;
        RECT 10.200 65.100 10.600 65.200 ;
        RECT 11.200 65.100 11.500 65.800 ;
        RECT 10.200 64.800 10.900 65.100 ;
        RECT 11.200 64.800 11.700 65.100 ;
        RECT 10.600 64.200 10.900 64.800 ;
        RECT 10.600 63.800 11.000 64.200 ;
        RECT 11.300 61.100 11.700 64.800 ;
        RECT 13.400 64.400 13.800 65.200 ;
        RECT 14.200 61.100 14.600 66.800 ;
        RECT 17.700 66.700 18.100 66.800 ;
        RECT 16.900 66.200 17.300 66.300 ;
        RECT 16.900 65.900 19.400 66.200 ;
        RECT 19.000 65.800 19.400 65.900 ;
        RECT 15.800 65.500 18.600 65.600 ;
        RECT 15.800 65.400 18.700 65.500 ;
        RECT 15.800 65.300 20.700 65.400 ;
        RECT 15.800 61.100 16.200 65.300 ;
        RECT 18.300 65.100 20.700 65.300 ;
        RECT 17.400 64.500 20.100 64.800 ;
        RECT 17.400 64.400 17.800 64.500 ;
        RECT 19.700 64.400 20.100 64.500 ;
        RECT 20.400 64.500 20.700 65.100 ;
        RECT 21.400 65.200 21.700 66.800 ;
        RECT 22.200 66.400 22.600 66.500 ;
        RECT 22.200 66.100 24.100 66.400 ;
        RECT 23.700 66.000 24.100 66.100 ;
        RECT 22.900 65.700 23.300 65.800 ;
        RECT 24.600 65.700 25.000 67.400 ;
        RECT 25.800 67.200 26.200 67.400 ;
        RECT 27.800 67.200 28.100 67.900 ;
        RECT 28.700 67.700 30.500 67.900 ;
        RECT 29.000 67.200 29.400 67.400 ;
        RECT 31.000 67.200 31.300 67.900 ;
        RECT 25.400 66.900 26.200 67.200 ;
        RECT 25.400 66.800 25.800 66.900 ;
        RECT 26.900 66.800 28.200 67.200 ;
        RECT 28.600 66.900 29.400 67.200 ;
        RECT 28.600 66.800 29.000 66.900 ;
        RECT 30.100 66.800 31.400 67.200 ;
        RECT 26.200 65.800 26.600 66.600 ;
        RECT 22.900 65.400 25.000 65.700 ;
        RECT 21.400 64.900 22.600 65.200 ;
        RECT 21.100 64.500 21.500 64.600 ;
        RECT 20.400 64.200 21.500 64.500 ;
        RECT 22.300 64.400 22.600 64.900 ;
        RECT 22.300 64.000 23.000 64.400 ;
        RECT 19.100 63.700 19.500 63.800 ;
        RECT 20.500 63.700 20.900 63.800 ;
        RECT 17.400 63.100 17.800 63.500 ;
        RECT 19.100 63.400 20.900 63.700 ;
        RECT 20.200 63.100 20.500 63.400 ;
        RECT 22.200 63.100 22.600 63.500 ;
        RECT 17.400 62.800 18.400 63.100 ;
        RECT 18.000 61.100 18.400 62.800 ;
        RECT 20.200 61.100 20.600 63.100 ;
        RECT 22.300 61.100 22.900 63.100 ;
        RECT 24.600 61.100 25.000 65.400 ;
        RECT 26.900 65.100 27.200 66.800 ;
        RECT 29.400 65.800 29.800 66.600 ;
        RECT 30.100 66.100 30.400 66.800 ;
        RECT 31.800 66.100 32.200 66.200 ;
        RECT 30.100 65.800 32.200 66.100 ;
        RECT 27.800 65.100 28.200 65.200 ;
        RECT 30.100 65.100 30.400 65.800 ;
        RECT 31.000 65.100 31.400 65.200 ;
        RECT 26.700 64.800 27.200 65.100 ;
        RECT 27.500 64.800 28.200 65.100 ;
        RECT 29.900 64.800 30.400 65.100 ;
        RECT 30.700 64.800 31.400 65.100 ;
        RECT 26.700 61.100 27.100 64.800 ;
        RECT 27.500 64.200 27.800 64.800 ;
        RECT 27.400 63.800 27.800 64.200 ;
        RECT 29.900 61.100 30.300 64.800 ;
        RECT 30.700 64.200 31.000 64.800 ;
        RECT 31.800 64.400 32.200 65.200 ;
        RECT 30.600 63.800 31.000 64.200 ;
        RECT 32.600 64.100 33.000 67.900 ;
        RECT 33.400 66.800 33.800 67.600 ;
        RECT 34.200 67.500 34.600 69.900 ;
        RECT 36.400 69.200 36.800 69.900 ;
        RECT 35.800 68.900 36.800 69.200 ;
        RECT 38.600 68.900 39.000 69.900 ;
        RECT 40.700 69.200 41.300 69.900 ;
        RECT 40.600 68.900 41.300 69.200 ;
        RECT 35.800 68.500 36.200 68.900 ;
        RECT 38.600 68.600 38.900 68.900 ;
        RECT 36.600 67.800 37.000 68.600 ;
        RECT 37.500 68.300 38.900 68.600 ;
        RECT 40.600 68.500 41.000 68.900 ;
        RECT 37.500 68.200 37.900 68.300 ;
        RECT 34.600 67.100 35.400 67.200 ;
        RECT 36.700 67.100 37.000 67.800 ;
        RECT 41.500 67.700 41.900 67.800 ;
        RECT 43.000 67.700 43.400 69.900 ;
        RECT 43.800 68.000 44.200 69.900 ;
        RECT 45.400 68.000 45.800 69.900 ;
        RECT 43.800 67.900 45.800 68.000 ;
        RECT 46.200 67.900 46.600 69.900 ;
        RECT 43.900 67.700 45.700 67.900 ;
        RECT 41.500 67.400 43.400 67.700 ;
        RECT 39.500 67.100 39.900 67.200 ;
        RECT 34.600 66.800 40.100 67.100 ;
        RECT 36.100 66.700 36.500 66.800 ;
        RECT 35.300 66.200 35.700 66.300 ;
        RECT 36.600 66.200 37.000 66.300 ;
        RECT 35.300 65.900 37.800 66.200 ;
        RECT 37.400 65.800 37.800 65.900 ;
        RECT 34.200 65.500 37.000 65.600 ;
        RECT 34.200 65.400 37.100 65.500 ;
        RECT 34.200 65.300 39.100 65.400 ;
        RECT 33.400 64.100 33.800 64.200 ;
        RECT 32.600 63.800 33.800 64.100 ;
        RECT 32.600 61.100 33.000 63.800 ;
        RECT 34.200 61.100 34.600 65.300 ;
        RECT 36.700 65.100 39.100 65.300 ;
        RECT 35.800 64.500 38.500 64.800 ;
        RECT 35.800 64.400 36.200 64.500 ;
        RECT 38.100 64.400 38.500 64.500 ;
        RECT 38.800 64.500 39.100 65.100 ;
        RECT 39.800 65.200 40.100 66.800 ;
        RECT 40.600 66.400 41.000 66.500 ;
        RECT 40.600 66.100 42.500 66.400 ;
        RECT 42.100 66.000 42.500 66.100 ;
        RECT 41.300 65.700 41.700 65.800 ;
        RECT 43.000 65.700 43.400 67.400 ;
        RECT 44.200 67.200 44.600 67.400 ;
        RECT 46.200 67.200 46.500 67.900 ;
        RECT 48.600 67.800 49.000 69.900 ;
        RECT 49.300 68.200 49.700 68.600 ;
        RECT 49.400 67.800 49.800 68.200 ;
        RECT 51.800 68.000 52.200 69.900 ;
        RECT 53.400 68.000 53.800 69.900 ;
        RECT 51.800 67.900 53.800 68.000 ;
        RECT 54.200 67.900 54.600 69.900 ;
        RECT 43.800 66.900 44.600 67.200 ;
        RECT 43.800 66.800 44.200 66.900 ;
        RECT 45.300 66.800 46.600 67.200 ;
        RECT 44.600 65.800 45.000 66.600 ;
        RECT 41.300 65.400 43.400 65.700 ;
        RECT 39.800 64.900 41.000 65.200 ;
        RECT 39.500 64.500 39.900 64.600 ;
        RECT 38.800 64.200 39.900 64.500 ;
        RECT 40.700 64.400 41.000 64.900 ;
        RECT 40.700 64.200 41.400 64.400 ;
        RECT 40.700 64.000 41.800 64.200 ;
        RECT 41.100 63.800 41.800 64.000 ;
        RECT 37.500 63.700 37.900 63.800 ;
        RECT 38.900 63.700 39.300 63.800 ;
        RECT 35.800 63.100 36.200 63.500 ;
        RECT 37.500 63.400 39.300 63.700 ;
        RECT 38.600 63.100 38.900 63.400 ;
        RECT 40.600 63.100 41.000 63.500 ;
        RECT 35.800 62.800 36.800 63.100 ;
        RECT 36.400 61.100 36.800 62.800 ;
        RECT 38.600 61.100 39.000 63.100 ;
        RECT 40.700 61.100 41.300 63.100 ;
        RECT 43.000 61.100 43.400 65.400 ;
        RECT 45.300 65.100 45.600 66.800 ;
        RECT 47.800 66.400 48.200 67.200 ;
        RECT 47.000 66.100 47.400 66.200 ;
        RECT 48.600 66.100 48.900 67.800 ;
        RECT 51.900 67.700 53.700 67.900 ;
        RECT 52.200 67.200 52.600 67.400 ;
        RECT 54.200 67.200 54.500 67.900 ;
        RECT 55.000 67.800 55.400 69.900 ;
        RECT 55.800 68.000 56.200 69.900 ;
        RECT 57.400 68.000 57.800 69.900 ;
        RECT 58.500 69.200 58.900 69.900 ;
        RECT 58.200 68.800 58.900 69.200 ;
        RECT 55.800 67.900 57.800 68.000 ;
        RECT 58.500 68.200 58.900 68.800 ;
        RECT 58.500 67.900 59.400 68.200 ;
        RECT 55.100 67.200 55.400 67.800 ;
        RECT 55.900 67.700 57.700 67.900 ;
        RECT 57.000 67.200 57.400 67.400 ;
        RECT 51.800 66.900 52.600 67.200 ;
        RECT 51.800 66.800 52.200 66.900 ;
        RECT 53.300 66.800 54.600 67.200 ;
        RECT 55.000 66.800 56.300 67.200 ;
        RECT 57.000 66.900 57.800 67.200 ;
        RECT 57.400 66.800 57.800 66.900 ;
        RECT 49.400 66.100 49.800 66.200 ;
        RECT 47.000 65.800 47.800 66.100 ;
        RECT 48.600 65.800 49.800 66.100 ;
        RECT 51.000 66.100 51.400 66.200 ;
        RECT 52.600 66.100 53.000 66.600 ;
        RECT 51.000 65.800 53.000 66.100 ;
        RECT 47.400 65.600 47.800 65.800 ;
        RECT 46.200 65.100 46.600 65.200 ;
        RECT 49.400 65.100 49.700 65.800 ;
        RECT 53.300 65.100 53.600 66.800 ;
        RECT 54.200 65.100 54.600 65.200 ;
        RECT 45.100 64.800 45.600 65.100 ;
        RECT 45.900 64.800 46.600 65.100 ;
        RECT 47.000 64.800 49.000 65.100 ;
        RECT 45.100 61.100 45.500 64.800 ;
        RECT 45.900 64.200 46.200 64.800 ;
        RECT 45.800 63.800 46.200 64.200 ;
        RECT 47.000 61.100 47.400 64.800 ;
        RECT 48.600 61.100 49.000 64.800 ;
        RECT 49.400 61.100 49.800 65.100 ;
        RECT 53.100 64.800 53.600 65.100 ;
        RECT 53.900 64.800 54.600 65.100 ;
        RECT 55.000 65.100 55.400 65.200 ;
        RECT 56.000 65.100 56.300 66.800 ;
        RECT 56.600 65.800 57.000 66.600 ;
        RECT 55.000 64.800 55.700 65.100 ;
        RECT 56.000 64.800 56.500 65.100 ;
        RECT 53.100 64.200 53.500 64.800 ;
        RECT 53.900 64.200 54.200 64.800 ;
        RECT 52.600 63.800 53.500 64.200 ;
        RECT 53.800 63.800 54.200 64.200 ;
        RECT 55.400 64.200 55.700 64.800 ;
        RECT 55.400 63.800 55.800 64.200 ;
        RECT 53.100 61.100 53.500 63.800 ;
        RECT 56.100 61.100 56.500 64.800 ;
        RECT 58.200 64.400 58.600 65.200 ;
        RECT 59.000 61.100 59.400 67.900 ;
        RECT 59.800 66.800 60.200 67.600 ;
        RECT 60.600 67.500 61.000 69.900 ;
        RECT 62.800 69.200 63.200 69.900 ;
        RECT 62.200 68.900 63.200 69.200 ;
        RECT 65.000 68.900 65.400 69.900 ;
        RECT 67.100 69.200 67.700 69.900 ;
        RECT 67.000 68.900 67.700 69.200 ;
        RECT 62.200 68.500 62.600 68.900 ;
        RECT 65.000 68.600 65.300 68.900 ;
        RECT 63.000 68.200 63.400 68.600 ;
        RECT 63.900 68.300 65.300 68.600 ;
        RECT 67.000 68.500 67.400 68.900 ;
        RECT 63.900 68.200 64.300 68.300 ;
        RECT 61.000 67.100 61.800 67.200 ;
        RECT 63.100 67.100 63.400 68.200 ;
        RECT 67.900 67.700 68.300 67.800 ;
        RECT 69.400 67.700 69.800 69.900 ;
        RECT 67.900 67.400 69.800 67.700 ;
        RECT 65.900 67.100 66.300 67.200 ;
        RECT 61.000 66.800 66.500 67.100 ;
        RECT 62.500 66.700 62.900 66.800 ;
        RECT 61.700 66.200 62.100 66.300 ;
        RECT 61.700 66.100 64.200 66.200 ;
        RECT 65.400 66.100 65.800 66.200 ;
        RECT 61.700 65.900 65.800 66.100 ;
        RECT 63.800 65.800 65.800 65.900 ;
        RECT 60.600 65.500 63.400 65.600 ;
        RECT 60.600 65.400 63.500 65.500 ;
        RECT 60.600 65.300 65.500 65.400 ;
        RECT 60.600 61.100 61.000 65.300 ;
        RECT 63.100 65.100 65.500 65.300 ;
        RECT 62.200 64.500 64.900 64.800 ;
        RECT 62.200 64.400 62.600 64.500 ;
        RECT 64.500 64.400 64.900 64.500 ;
        RECT 65.200 64.500 65.500 65.100 ;
        RECT 66.200 65.200 66.500 66.800 ;
        RECT 67.000 66.400 67.400 66.500 ;
        RECT 67.000 66.100 68.900 66.400 ;
        RECT 68.500 66.000 68.900 66.100 ;
        RECT 67.700 65.700 68.100 65.800 ;
        RECT 69.400 65.700 69.800 67.400 ;
        RECT 71.800 67.900 72.200 69.900 ;
        RECT 74.200 68.900 74.600 69.900 ;
        RECT 72.500 68.200 72.900 68.600 ;
        RECT 71.000 66.400 71.400 67.200 ;
        RECT 70.200 66.100 70.600 66.200 ;
        RECT 71.800 66.100 72.100 67.900 ;
        RECT 72.600 67.800 73.000 68.200 ;
        RECT 73.400 67.800 73.800 68.600 ;
        RECT 72.600 67.100 72.900 67.800 ;
        RECT 74.300 67.200 74.600 68.900 ;
        RECT 75.800 67.600 76.200 69.900 ;
        RECT 77.400 68.200 77.800 69.900 ;
        RECT 79.300 69.200 79.700 69.900 ;
        RECT 79.000 68.800 79.700 69.200 ;
        RECT 79.300 68.200 79.700 68.800 ;
        RECT 77.400 67.900 77.900 68.200 ;
        RECT 79.300 67.900 80.200 68.200 ;
        RECT 81.400 67.900 81.800 69.900 ;
        RECT 82.200 68.000 82.600 69.900 ;
        RECT 83.800 68.000 84.200 69.900 ;
        RECT 82.200 67.900 84.200 68.000 ;
        RECT 84.600 67.900 85.000 69.900 ;
        RECT 85.400 68.000 85.800 69.900 ;
        RECT 87.000 68.000 87.400 69.900 ;
        RECT 88.100 69.200 88.500 69.900 ;
        RECT 87.800 68.800 88.500 69.200 ;
        RECT 85.400 67.900 87.400 68.000 ;
        RECT 88.100 68.200 88.500 68.800 ;
        RECT 88.100 67.900 89.000 68.200 ;
        RECT 90.200 67.900 90.600 69.900 ;
        RECT 91.000 68.000 91.400 69.900 ;
        RECT 92.600 68.000 93.000 69.900 ;
        RECT 93.700 69.200 94.100 69.900 ;
        RECT 93.400 68.800 94.100 69.200 ;
        RECT 91.000 67.900 93.000 68.000 ;
        RECT 93.700 68.200 94.100 68.800 ;
        RECT 93.700 67.900 94.600 68.200 ;
        RECT 95.800 67.900 96.200 69.900 ;
        RECT 96.600 68.000 97.000 69.900 ;
        RECT 98.200 68.000 98.600 69.900 ;
        RECT 99.100 68.200 99.500 68.600 ;
        RECT 96.600 67.900 98.600 68.000 ;
        RECT 75.800 67.300 77.100 67.600 ;
        RECT 74.200 67.100 74.600 67.200 ;
        RECT 72.600 66.800 74.600 67.100 ;
        RECT 72.600 66.100 73.000 66.200 ;
        RECT 70.200 65.800 71.000 66.100 ;
        RECT 71.800 65.800 73.000 66.100 ;
        RECT 67.700 65.400 69.800 65.700 ;
        RECT 70.600 65.600 71.000 65.800 ;
        RECT 66.200 64.900 67.400 65.200 ;
        RECT 65.900 64.500 66.300 64.600 ;
        RECT 65.200 64.200 66.300 64.500 ;
        RECT 67.100 64.400 67.400 64.900 ;
        RECT 67.100 64.000 67.800 64.400 ;
        RECT 63.900 63.700 64.300 63.800 ;
        RECT 65.300 63.700 65.700 63.800 ;
        RECT 62.200 63.100 62.600 63.500 ;
        RECT 63.900 63.400 65.700 63.700 ;
        RECT 65.000 63.100 65.300 63.400 ;
        RECT 67.000 63.100 67.400 63.500 ;
        RECT 62.200 62.800 63.200 63.100 ;
        RECT 62.800 61.100 63.200 62.800 ;
        RECT 65.000 61.100 65.400 63.100 ;
        RECT 67.100 61.100 67.700 63.100 ;
        RECT 69.400 61.100 69.800 65.400 ;
        RECT 72.600 65.100 72.900 65.800 ;
        RECT 74.300 65.100 74.600 66.800 ;
        RECT 75.900 66.200 76.300 66.600 ;
        RECT 75.000 65.400 75.400 66.200 ;
        RECT 75.800 65.800 76.300 66.200 ;
        RECT 76.800 66.500 77.100 67.300 ;
        RECT 77.600 67.200 77.900 67.900 ;
        RECT 77.400 66.800 77.900 67.200 ;
        RECT 76.800 66.100 77.300 66.500 ;
        RECT 76.800 65.100 77.100 66.100 ;
        RECT 77.600 65.100 77.900 66.800 ;
        RECT 70.200 64.800 72.200 65.100 ;
        RECT 70.200 61.100 70.600 64.800 ;
        RECT 71.800 61.100 72.200 64.800 ;
        RECT 72.600 61.100 73.000 65.100 ;
        RECT 74.200 64.700 75.100 65.100 ;
        RECT 74.700 61.100 75.100 64.700 ;
        RECT 75.800 64.800 77.100 65.100 ;
        RECT 75.800 61.100 76.200 64.800 ;
        RECT 77.400 64.600 77.900 65.100 ;
        RECT 77.400 61.100 77.800 64.600 ;
        RECT 79.000 64.400 79.400 65.200 ;
        RECT 79.800 61.100 80.200 67.900 ;
        RECT 80.600 67.100 81.000 67.600 ;
        RECT 81.500 67.200 81.800 67.900 ;
        RECT 82.300 67.700 84.100 67.900 ;
        RECT 83.400 67.200 83.800 67.400 ;
        RECT 84.700 67.200 85.000 67.900 ;
        RECT 85.500 67.700 87.300 67.900 ;
        RECT 86.600 67.200 87.000 67.400 ;
        RECT 81.400 67.100 82.700 67.200 ;
        RECT 80.600 66.800 82.700 67.100 ;
        RECT 83.400 66.900 84.200 67.200 ;
        RECT 83.800 66.800 84.200 66.900 ;
        RECT 84.600 66.800 85.900 67.200 ;
        RECT 86.600 66.900 87.400 67.200 ;
        RECT 87.000 66.800 87.400 66.900 ;
        RECT 81.400 65.100 81.800 65.200 ;
        RECT 82.400 65.100 82.700 66.800 ;
        RECT 83.000 66.100 83.400 66.600 ;
        RECT 84.600 66.100 85.000 66.200 ;
        RECT 83.000 65.800 85.000 66.100 ;
        RECT 84.600 65.100 85.000 65.200 ;
        RECT 85.600 65.100 85.900 66.800 ;
        RECT 86.200 65.800 86.600 66.600 ;
        RECT 81.400 64.800 82.100 65.100 ;
        RECT 82.400 64.800 82.900 65.100 ;
        RECT 84.600 64.800 85.300 65.100 ;
        RECT 85.600 64.800 86.100 65.100 ;
        RECT 81.800 64.200 82.100 64.800 ;
        RECT 81.800 63.800 82.200 64.200 ;
        RECT 82.500 61.100 82.900 64.800 ;
        RECT 85.000 64.200 85.300 64.800 ;
        RECT 85.000 63.800 85.400 64.200 ;
        RECT 85.700 61.100 86.100 64.800 ;
        RECT 87.800 64.400 88.200 65.200 ;
        RECT 88.600 61.100 89.000 67.900 ;
        RECT 89.400 67.100 89.800 67.600 ;
        RECT 90.300 67.200 90.600 67.900 ;
        RECT 91.100 67.700 92.900 67.900 ;
        RECT 92.200 67.200 92.600 67.400 ;
        RECT 90.200 67.100 91.500 67.200 ;
        RECT 89.400 66.800 91.500 67.100 ;
        RECT 92.200 66.900 93.000 67.200 ;
        RECT 92.600 66.800 93.000 66.900 ;
        RECT 90.200 65.100 90.600 65.200 ;
        RECT 91.200 65.100 91.500 66.800 ;
        RECT 91.800 65.800 92.200 66.600 ;
        RECT 90.200 64.800 90.900 65.100 ;
        RECT 91.200 64.800 91.700 65.100 ;
        RECT 90.600 64.200 90.900 64.800 ;
        RECT 90.600 63.800 91.000 64.200 ;
        RECT 91.300 61.100 91.700 64.800 ;
        RECT 93.400 64.400 93.800 65.200 ;
        RECT 94.200 61.100 94.600 67.900 ;
        RECT 95.000 67.100 95.400 67.600 ;
        RECT 95.900 67.200 96.200 67.900 ;
        RECT 96.700 67.700 98.500 67.900 ;
        RECT 99.000 67.800 99.400 68.200 ;
        RECT 99.800 67.900 100.200 69.900 ;
        RECT 103.800 67.900 104.200 69.900 ;
        RECT 104.600 68.000 105.000 69.900 ;
        RECT 106.200 68.000 106.600 69.900 ;
        RECT 104.600 67.900 106.600 68.000 ;
        RECT 97.800 67.200 98.200 67.400 ;
        RECT 95.800 67.100 97.100 67.200 ;
        RECT 95.000 66.800 97.100 67.100 ;
        RECT 97.800 66.900 98.600 67.200 ;
        RECT 98.200 66.800 98.600 66.900 ;
        RECT 95.800 65.100 96.200 65.200 ;
        RECT 96.800 65.100 97.100 66.800 ;
        RECT 97.400 66.100 97.800 66.600 ;
        RECT 99.000 66.100 99.400 66.200 ;
        RECT 99.900 66.100 100.200 67.900 ;
        RECT 103.900 67.200 104.200 67.900 ;
        RECT 104.700 67.700 106.500 67.900 ;
        RECT 107.000 67.500 107.400 69.900 ;
        RECT 109.200 69.200 109.600 69.900 ;
        RECT 108.600 68.900 109.600 69.200 ;
        RECT 111.400 68.900 111.800 69.900 ;
        RECT 113.500 69.200 114.100 69.900 ;
        RECT 113.400 68.900 114.100 69.200 ;
        RECT 108.600 68.500 109.000 68.900 ;
        RECT 111.400 68.600 111.700 68.900 ;
        RECT 109.400 68.200 109.800 68.600 ;
        RECT 110.300 68.300 111.700 68.600 ;
        RECT 113.400 68.500 113.800 68.900 ;
        RECT 110.300 68.200 110.700 68.300 ;
        RECT 105.800 67.200 106.200 67.400 ;
        RECT 100.600 67.100 101.000 67.200 ;
        RECT 103.000 67.100 103.400 67.200 ;
        RECT 100.600 66.800 103.400 67.100 ;
        RECT 103.800 66.800 105.100 67.200 ;
        RECT 105.800 66.900 106.600 67.200 ;
        RECT 106.200 66.800 106.600 66.900 ;
        RECT 107.400 67.100 108.200 67.200 ;
        RECT 109.500 67.100 109.800 68.200 ;
        RECT 114.300 67.700 114.700 67.800 ;
        RECT 115.800 67.700 116.200 69.900 ;
        RECT 114.300 67.400 116.200 67.700 ;
        RECT 112.300 67.100 112.700 67.200 ;
        RECT 107.400 66.800 112.900 67.100 ;
        RECT 100.600 66.400 101.000 66.800 ;
        RECT 101.400 66.100 101.800 66.200 ;
        RECT 104.800 66.100 105.100 66.800 ;
        RECT 108.900 66.700 109.300 66.800 ;
        RECT 97.400 65.800 100.200 66.100 ;
        RECT 101.000 65.800 101.800 66.100 ;
        RECT 102.200 65.800 105.100 66.100 ;
        RECT 105.400 65.800 105.800 66.600 ;
        RECT 108.100 66.200 108.500 66.300 ;
        RECT 112.600 66.200 112.900 66.800 ;
        RECT 113.400 66.400 113.800 66.500 ;
        RECT 108.100 65.900 110.600 66.200 ;
        RECT 110.200 65.800 110.600 65.900 ;
        RECT 112.600 65.800 113.000 66.200 ;
        RECT 113.400 66.100 115.300 66.400 ;
        RECT 114.900 66.000 115.300 66.100 ;
        RECT 99.100 65.100 99.400 65.800 ;
        RECT 101.000 65.600 101.400 65.800 ;
        RECT 102.200 65.200 102.500 65.800 ;
        RECT 95.800 64.800 96.500 65.100 ;
        RECT 96.800 64.800 97.300 65.100 ;
        RECT 96.200 64.200 96.500 64.800 ;
        RECT 96.200 63.800 96.600 64.200 ;
        RECT 96.900 61.100 97.300 64.800 ;
        RECT 99.000 61.100 99.400 65.100 ;
        RECT 99.800 64.800 101.800 65.100 ;
        RECT 102.200 64.800 102.600 65.200 ;
        RECT 103.800 65.100 104.200 65.200 ;
        RECT 104.800 65.100 105.100 65.800 ;
        RECT 107.000 65.500 109.800 65.600 ;
        RECT 107.000 65.400 109.900 65.500 ;
        RECT 107.000 65.300 111.900 65.400 ;
        RECT 103.800 64.800 104.500 65.100 ;
        RECT 104.800 64.800 105.300 65.100 ;
        RECT 99.800 61.100 100.200 64.800 ;
        RECT 101.400 61.100 101.800 64.800 ;
        RECT 104.200 64.200 104.500 64.800 ;
        RECT 104.200 63.800 104.600 64.200 ;
        RECT 104.900 61.100 105.300 64.800 ;
        RECT 107.000 61.100 107.400 65.300 ;
        RECT 109.500 65.100 111.900 65.300 ;
        RECT 108.600 64.500 111.300 64.800 ;
        RECT 108.600 64.400 109.000 64.500 ;
        RECT 110.900 64.400 111.300 64.500 ;
        RECT 111.600 64.500 111.900 65.100 ;
        RECT 112.600 65.200 112.900 65.800 ;
        RECT 114.100 65.700 114.500 65.800 ;
        RECT 115.800 65.700 116.200 67.400 ;
        RECT 118.200 67.800 118.600 69.900 ;
        RECT 118.900 68.200 119.300 68.600 ;
        RECT 119.000 67.800 119.400 68.200 ;
        RECT 117.400 66.400 117.800 67.200 ;
        RECT 116.600 66.100 117.000 66.200 ;
        RECT 118.200 66.100 118.500 67.800 ;
        RECT 119.800 67.700 120.200 69.900 ;
        RECT 121.900 69.200 122.500 69.900 ;
        RECT 121.900 68.900 122.600 69.200 ;
        RECT 124.200 68.900 124.600 69.900 ;
        RECT 126.400 69.200 126.800 69.900 ;
        RECT 126.400 68.900 127.400 69.200 ;
        RECT 122.200 68.500 122.600 68.900 ;
        RECT 124.300 68.600 124.600 68.900 ;
        RECT 124.300 68.300 125.700 68.600 ;
        RECT 125.300 68.200 125.700 68.300 ;
        RECT 126.200 68.200 126.600 68.600 ;
        RECT 127.000 68.500 127.400 68.900 ;
        RECT 123.000 68.100 123.400 68.200 ;
        RECT 121.400 67.800 123.400 68.100 ;
        RECT 121.300 67.700 121.800 67.800 ;
        RECT 119.800 67.400 121.800 67.700 ;
        RECT 119.000 67.100 119.400 67.200 ;
        RECT 119.800 67.100 120.200 67.400 ;
        RECT 123.300 67.100 123.700 67.200 ;
        RECT 126.200 67.100 126.500 68.200 ;
        RECT 128.600 67.500 129.000 69.900 ;
        RECT 129.500 68.200 129.900 68.600 ;
        RECT 129.400 67.800 129.800 68.200 ;
        RECT 130.200 67.900 130.600 69.900 ;
        RECT 133.900 68.200 134.300 69.900 ;
        RECT 127.800 67.100 128.600 67.200 ;
        RECT 119.000 66.800 120.200 67.100 ;
        RECT 119.000 66.100 119.400 66.200 ;
        RECT 116.600 65.800 117.400 66.100 ;
        RECT 118.200 65.800 119.400 66.100 ;
        RECT 114.100 65.400 116.200 65.700 ;
        RECT 117.000 65.600 117.400 65.800 ;
        RECT 112.600 64.900 113.800 65.200 ;
        RECT 112.300 64.500 112.700 64.600 ;
        RECT 111.600 64.200 112.700 64.500 ;
        RECT 113.500 64.400 113.800 64.900 ;
        RECT 113.500 64.000 114.200 64.400 ;
        RECT 110.300 63.700 110.700 63.800 ;
        RECT 111.700 63.700 112.100 63.800 ;
        RECT 108.600 63.100 109.000 63.500 ;
        RECT 110.300 63.400 112.100 63.700 ;
        RECT 111.400 63.100 111.700 63.400 ;
        RECT 113.400 63.100 113.800 63.500 ;
        RECT 108.600 62.800 109.600 63.100 ;
        RECT 109.200 61.100 109.600 62.800 ;
        RECT 111.400 61.100 111.800 63.100 ;
        RECT 113.500 61.100 114.100 63.100 ;
        RECT 115.800 61.100 116.200 65.400 ;
        RECT 119.000 65.100 119.300 65.800 ;
        RECT 119.800 65.700 120.200 66.800 ;
        RECT 123.100 66.800 128.600 67.100 ;
        RECT 122.200 66.400 122.600 66.500 ;
        RECT 120.700 66.100 122.600 66.400 ;
        RECT 120.700 66.000 121.100 66.100 ;
        RECT 121.500 65.700 121.900 65.800 ;
        RECT 119.800 65.400 121.900 65.700 ;
        RECT 116.600 64.800 118.600 65.100 ;
        RECT 116.600 61.100 117.000 64.800 ;
        RECT 118.200 61.100 118.600 64.800 ;
        RECT 119.000 61.100 119.400 65.100 ;
        RECT 119.800 61.100 120.200 65.400 ;
        RECT 123.100 65.200 123.400 66.800 ;
        RECT 126.700 66.700 127.100 66.800 ;
        RECT 126.200 66.200 126.600 66.300 ;
        RECT 127.500 66.200 127.900 66.300 ;
        RECT 130.300 66.200 130.600 67.900 ;
        RECT 133.400 67.900 134.300 68.200 ;
        RECT 131.000 66.400 131.400 67.200 ;
        RECT 132.600 66.800 133.000 67.600 ;
        RECT 125.400 65.900 127.900 66.200 ;
        RECT 129.400 66.100 129.800 66.200 ;
        RECT 130.200 66.100 130.600 66.200 ;
        RECT 131.800 66.100 132.200 66.200 ;
        RECT 132.600 66.100 133.000 66.200 ;
        RECT 125.400 65.800 125.800 65.900 ;
        RECT 129.400 65.800 130.600 66.100 ;
        RECT 131.400 65.800 133.000 66.100 ;
        RECT 133.400 66.100 133.800 67.900 ;
        RECT 135.000 67.800 135.400 69.900 ;
        RECT 135.800 68.000 136.200 69.900 ;
        RECT 137.400 68.000 137.800 69.900 ;
        RECT 135.800 67.900 137.800 68.000 ;
        RECT 139.800 67.900 140.200 69.900 ;
        RECT 140.500 68.200 140.900 68.600 ;
        RECT 135.100 67.200 135.400 67.800 ;
        RECT 135.900 67.700 137.700 67.900 ;
        RECT 137.000 67.200 137.400 67.400 ;
        RECT 135.000 66.800 136.300 67.200 ;
        RECT 137.000 66.900 137.800 67.200 ;
        RECT 137.400 66.800 137.800 66.900 ;
        RECT 133.400 65.800 135.300 66.100 ;
        RECT 126.200 65.500 129.000 65.600 ;
        RECT 126.100 65.400 129.000 65.500 ;
        RECT 122.200 64.900 123.400 65.200 ;
        RECT 124.100 65.300 129.000 65.400 ;
        RECT 124.100 65.100 126.500 65.300 ;
        RECT 122.200 64.400 122.500 64.900 ;
        RECT 121.800 64.000 122.500 64.400 ;
        RECT 123.300 64.500 123.700 64.600 ;
        RECT 124.100 64.500 124.400 65.100 ;
        RECT 123.300 64.200 124.400 64.500 ;
        RECT 124.700 64.500 127.400 64.800 ;
        RECT 124.700 64.400 125.100 64.500 ;
        RECT 127.000 64.400 127.400 64.500 ;
        RECT 123.900 63.700 124.300 63.800 ;
        RECT 125.300 63.700 125.700 63.800 ;
        RECT 122.200 63.100 122.600 63.500 ;
        RECT 123.900 63.400 125.700 63.700 ;
        RECT 124.300 63.100 124.600 63.400 ;
        RECT 127.000 63.100 127.400 63.500 ;
        RECT 121.900 61.100 122.500 63.100 ;
        RECT 124.200 61.100 124.600 63.100 ;
        RECT 126.400 62.800 127.400 63.100 ;
        RECT 126.400 61.100 126.800 62.800 ;
        RECT 128.600 61.100 129.000 65.300 ;
        RECT 129.500 65.100 129.800 65.800 ;
        RECT 131.400 65.600 131.800 65.800 ;
        RECT 129.400 61.100 129.800 65.100 ;
        RECT 130.200 64.800 132.200 65.100 ;
        RECT 130.200 61.100 130.600 64.800 ;
        RECT 131.800 61.100 132.200 64.800 ;
        RECT 133.400 61.100 133.800 65.800 ;
        RECT 135.000 65.200 135.300 65.800 ;
        RECT 134.200 64.400 134.600 65.200 ;
        RECT 135.000 65.100 135.400 65.200 ;
        RECT 136.000 65.100 136.300 66.800 ;
        RECT 136.600 65.800 137.000 66.600 ;
        RECT 139.000 66.400 139.400 67.200 ;
        RECT 138.200 66.100 138.600 66.200 ;
        RECT 139.800 66.100 140.100 67.900 ;
        RECT 140.600 67.800 141.000 68.200 ;
        RECT 141.400 67.600 141.800 69.900 ;
        RECT 143.000 68.200 143.400 69.900 ;
        RECT 143.000 67.900 143.500 68.200 ;
        RECT 141.400 67.300 142.700 67.600 ;
        RECT 141.500 66.200 141.900 66.600 ;
        RECT 140.600 66.100 141.000 66.200 ;
        RECT 138.200 65.800 139.000 66.100 ;
        RECT 139.800 65.800 141.000 66.100 ;
        RECT 141.400 65.800 141.900 66.200 ;
        RECT 142.400 66.500 142.700 67.300 ;
        RECT 143.200 67.200 143.500 67.900 ;
        RECT 144.600 67.800 145.000 69.900 ;
        RECT 145.400 68.000 145.800 69.900 ;
        RECT 147.000 68.000 147.400 69.900 ;
        RECT 145.400 67.900 147.400 68.000 ;
        RECT 149.400 67.900 149.800 69.900 ;
        RECT 150.100 68.200 150.500 68.600 ;
        RECT 144.700 67.200 145.000 67.800 ;
        RECT 145.500 67.700 147.300 67.900 ;
        RECT 146.600 67.200 147.000 67.400 ;
        RECT 143.000 67.100 143.500 67.200 ;
        RECT 143.000 66.800 144.100 67.100 ;
        RECT 144.600 66.800 145.900 67.200 ;
        RECT 146.600 66.900 147.400 67.200 ;
        RECT 147.000 66.800 147.400 66.900 ;
        RECT 147.800 67.100 148.200 67.200 ;
        RECT 148.600 67.100 149.000 67.200 ;
        RECT 147.800 66.800 149.000 67.100 ;
        RECT 142.400 66.100 142.900 66.500 ;
        RECT 138.600 65.600 139.000 65.800 ;
        RECT 140.600 65.100 140.900 65.800 ;
        RECT 142.400 65.100 142.700 66.100 ;
        RECT 143.200 65.100 143.500 66.800 ;
        RECT 143.800 66.100 144.100 66.800 ;
        RECT 144.600 66.100 145.000 66.200 ;
        RECT 143.800 65.800 145.000 66.100 ;
        RECT 135.000 64.800 135.700 65.100 ;
        RECT 136.000 64.800 136.500 65.100 ;
        RECT 135.400 64.200 135.700 64.800 ;
        RECT 135.400 63.800 135.800 64.200 ;
        RECT 136.100 61.100 136.500 64.800 ;
        RECT 138.200 64.800 140.200 65.100 ;
        RECT 138.200 61.100 138.600 64.800 ;
        RECT 139.800 61.100 140.200 64.800 ;
        RECT 140.600 61.100 141.000 65.100 ;
        RECT 141.400 64.800 142.700 65.100 ;
        RECT 141.400 61.100 141.800 64.800 ;
        RECT 143.000 64.600 143.500 65.100 ;
        RECT 144.600 65.200 144.900 65.800 ;
        RECT 144.600 65.100 145.000 65.200 ;
        RECT 145.600 65.100 145.900 66.800 ;
        RECT 146.200 65.800 146.600 66.600 ;
        RECT 148.600 66.400 149.000 66.800 ;
        RECT 147.800 66.100 148.200 66.200 ;
        RECT 149.400 66.100 149.700 67.900 ;
        RECT 150.200 67.800 150.600 68.200 ;
        RECT 151.000 68.000 151.400 69.900 ;
        RECT 152.600 68.000 153.000 69.900 ;
        RECT 151.000 67.900 153.000 68.000 ;
        RECT 151.100 67.700 152.900 67.900 ;
        RECT 153.400 67.800 153.800 69.900 ;
        RECT 151.400 67.200 151.800 67.400 ;
        RECT 153.400 67.200 153.700 67.800 ;
        RECT 155.800 67.500 156.200 69.900 ;
        RECT 158.000 69.200 158.400 69.900 ;
        RECT 157.400 68.900 158.400 69.200 ;
        RECT 160.200 68.900 160.600 69.900 ;
        RECT 162.300 69.200 162.900 69.900 ;
        RECT 162.200 68.900 162.900 69.200 ;
        RECT 157.400 68.500 157.800 68.900 ;
        RECT 160.200 68.600 160.500 68.900 ;
        RECT 158.200 68.200 158.600 68.600 ;
        RECT 159.100 68.300 160.500 68.600 ;
        RECT 162.200 68.500 162.600 68.900 ;
        RECT 159.100 68.200 159.500 68.300 ;
        RECT 151.000 66.900 151.800 67.200 ;
        RECT 151.000 66.800 151.400 66.900 ;
        RECT 152.500 66.800 153.800 67.200 ;
        RECT 156.200 67.100 157.000 67.200 ;
        RECT 158.300 67.100 158.600 68.200 ;
        RECT 163.000 67.800 163.400 68.200 ;
        RECT 163.000 67.700 163.500 67.800 ;
        RECT 164.600 67.700 165.000 69.900 ;
        RECT 163.000 67.400 165.000 67.700 ;
        RECT 161.100 67.100 161.500 67.200 ;
        RECT 156.200 66.800 161.700 67.100 ;
        RECT 150.200 66.100 150.600 66.200 ;
        RECT 147.800 65.800 148.600 66.100 ;
        RECT 149.400 65.800 150.600 66.100 ;
        RECT 151.800 65.800 152.200 66.600 ;
        RECT 148.200 65.600 148.600 65.800 ;
        RECT 150.200 65.100 150.500 65.800 ;
        RECT 152.500 65.100 152.800 66.800 ;
        RECT 157.700 66.700 158.100 66.800 ;
        RECT 156.900 66.200 157.300 66.300 ;
        RECT 158.200 66.200 158.600 66.300 ;
        RECT 156.900 65.900 159.400 66.200 ;
        RECT 159.000 65.800 159.400 65.900 ;
        RECT 155.800 65.500 158.600 65.600 ;
        RECT 155.800 65.400 158.700 65.500 ;
        RECT 155.800 65.300 160.700 65.400 ;
        RECT 153.400 65.100 153.800 65.200 ;
        RECT 154.200 65.100 154.600 65.200 ;
        RECT 144.600 64.800 145.300 65.100 ;
        RECT 145.600 64.800 146.100 65.100 ;
        RECT 143.000 61.100 143.400 64.600 ;
        RECT 145.000 64.200 145.300 64.800 ;
        RECT 145.000 63.800 145.400 64.200 ;
        RECT 145.700 61.100 146.100 64.800 ;
        RECT 147.800 64.800 149.800 65.100 ;
        RECT 147.800 61.100 148.200 64.800 ;
        RECT 149.400 61.100 149.800 64.800 ;
        RECT 150.200 61.100 150.600 65.100 ;
        RECT 152.300 64.800 152.800 65.100 ;
        RECT 153.100 64.800 154.600 65.100 ;
        RECT 152.300 61.100 152.700 64.800 ;
        RECT 153.100 64.200 153.400 64.800 ;
        RECT 153.000 63.800 153.400 64.200 ;
        RECT 155.800 61.100 156.200 65.300 ;
        RECT 158.300 65.100 160.700 65.300 ;
        RECT 157.400 64.500 160.100 64.800 ;
        RECT 157.400 64.400 157.800 64.500 ;
        RECT 159.700 64.400 160.100 64.500 ;
        RECT 160.400 64.500 160.700 65.100 ;
        RECT 161.400 65.200 161.700 66.800 ;
        RECT 162.200 66.400 162.600 66.500 ;
        RECT 162.200 66.100 164.100 66.400 ;
        RECT 163.700 66.000 164.100 66.100 ;
        RECT 162.900 65.700 163.300 65.800 ;
        RECT 164.600 65.700 165.000 67.400 ;
        RECT 165.400 68.500 165.800 69.500 ;
        RECT 165.400 67.400 165.700 68.500 ;
        RECT 167.500 68.000 167.900 69.500 ;
        RECT 167.500 67.700 168.300 68.000 ;
        RECT 167.900 67.500 168.300 67.700 ;
        RECT 165.400 67.100 167.500 67.400 ;
        RECT 167.000 66.900 167.500 67.100 ;
        RECT 168.000 67.200 168.300 67.500 ;
        RECT 165.400 65.800 165.800 66.600 ;
        RECT 166.200 65.800 166.600 66.600 ;
        RECT 167.000 66.500 167.700 66.900 ;
        RECT 168.000 66.800 169.000 67.200 ;
        RECT 170.200 67.100 170.600 69.900 ;
        RECT 171.000 68.100 171.400 68.600 ;
        RECT 171.800 68.100 172.200 69.900 ;
        RECT 173.900 69.200 174.500 69.900 ;
        RECT 173.900 68.900 174.600 69.200 ;
        RECT 176.200 68.900 176.600 69.900 ;
        RECT 178.400 69.200 178.800 69.900 ;
        RECT 178.400 68.900 179.400 69.200 ;
        RECT 174.200 68.500 174.600 68.900 ;
        RECT 176.300 68.600 176.600 68.900 ;
        RECT 176.300 68.300 177.700 68.600 ;
        RECT 177.300 68.200 177.700 68.300 ;
        RECT 178.200 68.200 178.600 68.600 ;
        RECT 179.000 68.500 179.400 68.900 ;
        RECT 171.000 67.800 172.200 68.100 ;
        RECT 169.400 66.800 170.600 67.100 ;
        RECT 162.900 65.400 165.000 65.700 ;
        RECT 167.000 65.500 167.300 66.500 ;
        RECT 161.400 64.900 162.600 65.200 ;
        RECT 161.100 64.500 161.500 64.600 ;
        RECT 160.400 64.200 161.500 64.500 ;
        RECT 162.300 64.400 162.600 64.900 ;
        RECT 162.300 64.000 163.000 64.400 ;
        RECT 159.100 63.700 159.500 63.800 ;
        RECT 160.500 63.700 160.900 63.800 ;
        RECT 157.400 63.100 157.800 63.500 ;
        RECT 159.100 63.400 160.900 63.700 ;
        RECT 160.200 63.100 160.500 63.400 ;
        RECT 162.200 63.100 162.600 63.500 ;
        RECT 157.400 62.800 158.400 63.100 ;
        RECT 158.000 61.100 158.400 62.800 ;
        RECT 160.200 61.100 160.600 63.100 ;
        RECT 162.300 61.100 162.900 63.100 ;
        RECT 164.600 61.100 165.000 65.400 ;
        RECT 165.400 65.200 167.300 65.500 ;
        RECT 168.000 65.200 168.300 66.800 ;
        RECT 169.400 66.200 169.700 66.800 ;
        RECT 168.600 65.400 169.000 66.200 ;
        RECT 169.400 65.800 169.800 66.200 ;
        RECT 165.400 63.500 165.700 65.200 ;
        RECT 167.800 64.900 168.300 65.200 ;
        RECT 167.500 64.600 168.300 64.900 ;
        RECT 165.400 61.500 165.800 63.500 ;
        RECT 167.500 61.100 167.900 64.600 ;
        RECT 170.200 61.100 170.600 66.800 ;
        RECT 171.800 67.700 172.200 67.800 ;
        RECT 173.300 67.700 173.700 67.800 ;
        RECT 171.800 67.400 173.700 67.700 ;
        RECT 171.800 65.700 172.200 67.400 ;
        RECT 175.300 67.100 175.700 67.200 ;
        RECT 178.200 67.100 178.500 68.200 ;
        RECT 180.600 67.500 181.000 69.900 ;
        RECT 183.300 68.000 183.700 69.500 ;
        RECT 185.400 68.500 185.800 69.500 ;
        RECT 182.900 67.700 183.700 68.000 ;
        RECT 182.900 67.500 183.300 67.700 ;
        RECT 182.900 67.200 183.200 67.500 ;
        RECT 185.500 67.400 185.800 68.500 ;
        RECT 179.800 67.100 180.600 67.200 ;
        RECT 181.400 67.100 181.800 67.200 ;
        RECT 175.100 66.800 181.800 67.100 ;
        RECT 182.200 66.800 183.200 67.200 ;
        RECT 183.700 67.100 185.800 67.400 ;
        RECT 187.800 67.800 188.200 69.900 ;
        RECT 188.500 68.200 188.900 68.600 ;
        RECT 188.600 68.100 189.000 68.200 ;
        RECT 189.400 68.100 189.800 69.900 ;
        RECT 188.600 67.800 189.800 68.100 ;
        RECT 190.200 68.000 190.600 69.900 ;
        RECT 191.800 68.000 192.200 69.900 ;
        RECT 190.200 67.900 192.200 68.000 ;
        RECT 183.700 66.900 184.200 67.100 ;
        RECT 174.200 66.400 174.600 66.500 ;
        RECT 172.700 66.100 174.600 66.400 ;
        RECT 175.100 66.200 175.400 66.800 ;
        RECT 178.700 66.700 179.100 66.800 ;
        RECT 179.500 66.200 179.900 66.300 ;
        RECT 172.700 66.000 173.100 66.100 ;
        RECT 175.000 65.800 175.400 66.200 ;
        RECT 175.800 66.100 176.200 66.200 ;
        RECT 177.400 66.100 179.900 66.200 ;
        RECT 175.800 65.900 179.900 66.100 ;
        RECT 175.800 65.800 177.800 65.900 ;
        RECT 173.500 65.700 173.900 65.800 ;
        RECT 171.800 65.400 173.900 65.700 ;
        RECT 171.800 61.100 172.200 65.400 ;
        RECT 175.100 65.200 175.400 65.800 ;
        RECT 178.200 65.500 181.000 65.600 ;
        RECT 178.100 65.400 181.000 65.500 ;
        RECT 182.200 65.400 182.600 66.200 ;
        RECT 174.200 64.900 175.400 65.200 ;
        RECT 176.100 65.300 181.000 65.400 ;
        RECT 176.100 65.100 178.500 65.300 ;
        RECT 174.200 64.400 174.500 64.900 ;
        RECT 173.800 64.000 174.500 64.400 ;
        RECT 175.300 64.500 175.700 64.600 ;
        RECT 176.100 64.500 176.400 65.100 ;
        RECT 175.300 64.200 176.400 64.500 ;
        RECT 176.700 64.500 179.400 64.800 ;
        RECT 176.700 64.400 177.100 64.500 ;
        RECT 179.000 64.400 179.400 64.500 ;
        RECT 175.900 63.700 176.300 63.800 ;
        RECT 177.300 63.700 177.700 63.800 ;
        RECT 174.200 63.100 174.600 63.500 ;
        RECT 175.900 63.400 177.700 63.700 ;
        RECT 176.300 63.100 176.600 63.400 ;
        RECT 179.000 63.100 179.400 63.500 ;
        RECT 173.900 61.100 174.500 63.100 ;
        RECT 176.200 61.100 176.600 63.100 ;
        RECT 178.400 62.800 179.400 63.100 ;
        RECT 178.400 61.100 178.800 62.800 ;
        RECT 180.600 61.100 181.000 65.300 ;
        RECT 182.900 64.900 183.200 66.800 ;
        RECT 183.500 66.500 184.200 66.900 ;
        RECT 183.900 65.500 184.200 66.500 ;
        RECT 184.600 65.800 185.000 66.600 ;
        RECT 185.400 65.800 185.800 66.600 ;
        RECT 187.000 66.400 187.400 67.200 ;
        RECT 186.200 66.100 186.600 66.200 ;
        RECT 187.800 66.100 188.100 67.800 ;
        RECT 189.500 67.200 189.800 67.800 ;
        RECT 190.300 67.700 192.100 67.900 ;
        RECT 191.400 67.200 191.800 67.400 ;
        RECT 189.400 66.800 190.700 67.200 ;
        RECT 191.400 66.900 192.200 67.200 ;
        RECT 191.800 66.800 192.200 66.900 ;
        RECT 188.600 66.100 189.000 66.200 ;
        RECT 186.200 65.800 187.000 66.100 ;
        RECT 187.800 65.800 189.000 66.100 ;
        RECT 186.600 65.600 187.000 65.800 ;
        RECT 183.900 65.200 185.800 65.500 ;
        RECT 182.900 64.600 183.700 64.900 ;
        RECT 183.300 62.200 183.700 64.600 ;
        RECT 185.500 63.500 185.800 65.200 ;
        RECT 188.600 65.100 188.900 65.800 ;
        RECT 189.400 65.100 189.800 65.200 ;
        RECT 190.400 65.100 190.700 66.800 ;
        RECT 191.000 65.800 191.400 66.600 ;
        RECT 191.800 66.100 192.200 66.200 ;
        RECT 193.400 66.100 193.800 69.900 ;
        RECT 195.000 67.900 195.400 69.900 ;
        RECT 195.800 68.000 196.200 69.900 ;
        RECT 197.400 68.000 197.800 69.900 ;
        RECT 199.000 68.800 199.400 69.900 ;
        RECT 195.800 67.900 197.800 68.000 ;
        RECT 195.100 67.200 195.400 67.900 ;
        RECT 195.900 67.700 197.700 67.900 ;
        RECT 198.200 67.800 198.600 68.600 ;
        RECT 197.000 67.200 197.400 67.400 ;
        RECT 199.100 67.200 199.400 68.800 ;
        RECT 200.700 68.200 201.100 68.600 ;
        RECT 200.600 67.800 201.000 68.200 ;
        RECT 201.400 67.900 201.800 69.900 ;
        RECT 195.000 66.800 196.300 67.200 ;
        RECT 197.000 66.900 197.800 67.200 ;
        RECT 197.400 66.800 197.800 66.900 ;
        RECT 199.000 66.800 199.400 67.200 ;
        RECT 191.800 65.800 193.800 66.100 ;
        RECT 183.000 61.800 183.700 62.200 ;
        RECT 183.300 61.100 183.700 61.800 ;
        RECT 185.400 61.500 185.800 63.500 ;
        RECT 186.200 64.800 188.200 65.100 ;
        RECT 186.200 61.100 186.600 64.800 ;
        RECT 187.800 61.100 188.200 64.800 ;
        RECT 188.600 61.100 189.000 65.100 ;
        RECT 189.400 64.800 190.100 65.100 ;
        RECT 190.400 64.800 190.900 65.100 ;
        RECT 189.800 64.200 190.100 64.800 ;
        RECT 189.800 63.800 190.200 64.200 ;
        RECT 190.500 61.100 190.900 64.800 ;
        RECT 193.400 61.100 193.800 65.800 ;
        RECT 195.000 65.100 195.400 65.200 ;
        RECT 196.000 65.100 196.300 66.800 ;
        RECT 196.600 65.800 197.000 66.600 ;
        RECT 199.100 65.100 199.400 66.800 ;
        RECT 199.800 65.400 200.200 66.200 ;
        RECT 200.600 66.100 201.000 66.200 ;
        RECT 201.500 66.100 201.800 67.900 ;
        RECT 202.200 66.400 202.600 67.200 ;
        RECT 203.000 66.100 203.400 66.200 ;
        RECT 200.600 65.800 201.800 66.100 ;
        RECT 202.600 65.800 203.400 66.100 ;
        RECT 200.700 65.100 201.000 65.800 ;
        RECT 202.600 65.600 203.000 65.800 ;
        RECT 195.000 64.800 195.700 65.100 ;
        RECT 196.000 64.800 196.500 65.100 ;
        RECT 195.400 64.200 195.700 64.800 ;
        RECT 195.400 63.800 195.800 64.200 ;
        RECT 196.100 61.100 196.500 64.800 ;
        RECT 199.000 64.700 199.900 65.100 ;
        RECT 199.500 61.100 199.900 64.700 ;
        RECT 200.600 61.100 201.000 65.100 ;
        RECT 201.400 64.800 203.400 65.100 ;
        RECT 201.400 61.100 201.800 64.800 ;
        RECT 203.000 61.100 203.400 64.800 ;
        RECT 0.600 55.700 1.000 59.900 ;
        RECT 2.800 58.200 3.200 59.900 ;
        RECT 2.200 57.900 3.200 58.200 ;
        RECT 5.000 57.900 5.400 59.900 ;
        RECT 7.100 57.900 7.700 59.900 ;
        RECT 2.200 57.500 2.600 57.900 ;
        RECT 5.000 57.600 5.300 57.900 ;
        RECT 3.900 57.300 5.700 57.600 ;
        RECT 7.000 57.500 7.400 57.900 ;
        RECT 3.900 57.200 4.300 57.300 ;
        RECT 5.300 57.200 5.700 57.300 ;
        RECT 2.200 56.500 2.600 56.600 ;
        RECT 4.500 56.500 4.900 56.600 ;
        RECT 2.200 56.200 4.900 56.500 ;
        RECT 5.200 56.500 6.300 56.800 ;
        RECT 5.200 55.900 5.500 56.500 ;
        RECT 5.900 56.400 6.300 56.500 ;
        RECT 7.100 56.600 7.800 57.000 ;
        RECT 7.100 56.100 7.400 56.600 ;
        RECT 3.100 55.700 5.500 55.900 ;
        RECT 0.600 55.600 5.500 55.700 ;
        RECT 6.200 55.800 7.400 56.100 ;
        RECT 0.600 55.500 3.500 55.600 ;
        RECT 0.600 55.400 3.400 55.500 ;
        RECT 3.800 55.100 4.200 55.200 ;
        RECT 1.700 54.800 4.200 55.100 ;
        RECT 1.700 54.700 2.100 54.800 ;
        RECT 2.500 54.200 2.900 54.300 ;
        RECT 6.200 54.200 6.500 55.800 ;
        RECT 9.400 55.600 9.800 59.900 ;
        RECT 7.700 55.300 9.800 55.600 ;
        RECT 10.200 55.700 10.600 59.900 ;
        RECT 12.400 58.200 12.800 59.900 ;
        RECT 11.800 57.900 12.800 58.200 ;
        RECT 14.600 57.900 15.000 59.900 ;
        RECT 16.700 57.900 17.300 59.900 ;
        RECT 11.800 57.500 12.200 57.900 ;
        RECT 14.600 57.600 14.900 57.900 ;
        RECT 13.500 57.300 15.300 57.600 ;
        RECT 16.600 57.500 17.000 57.900 ;
        RECT 13.500 57.200 13.900 57.300 ;
        RECT 14.900 57.200 15.300 57.300 ;
        RECT 11.800 56.500 12.200 56.600 ;
        RECT 14.100 56.500 14.500 56.600 ;
        RECT 11.800 56.200 14.500 56.500 ;
        RECT 14.800 56.500 15.900 56.800 ;
        RECT 14.800 55.900 15.100 56.500 ;
        RECT 15.500 56.400 15.900 56.500 ;
        RECT 16.700 56.600 17.400 57.000 ;
        RECT 16.700 56.100 17.000 56.600 ;
        RECT 12.700 55.700 15.100 55.900 ;
        RECT 10.200 55.600 15.100 55.700 ;
        RECT 15.800 55.800 17.000 56.100 ;
        RECT 10.200 55.500 13.100 55.600 ;
        RECT 10.200 55.400 13.000 55.500 ;
        RECT 7.700 55.200 8.100 55.300 ;
        RECT 8.500 54.900 8.900 55.000 ;
        RECT 7.000 54.600 8.900 54.900 ;
        RECT 7.000 54.500 7.400 54.600 ;
        RECT 1.000 53.900 6.500 54.200 ;
        RECT 1.000 53.800 1.800 53.900 ;
        RECT 0.600 51.100 1.000 53.500 ;
        RECT 3.100 53.200 3.400 53.900 ;
        RECT 5.900 53.800 6.300 53.900 ;
        RECT 9.400 53.600 9.800 55.300 ;
        RECT 13.400 55.100 13.800 55.200 ;
        RECT 14.200 55.100 14.600 55.200 ;
        RECT 11.300 54.800 14.600 55.100 ;
        RECT 11.300 54.700 11.700 54.800 ;
        RECT 12.100 54.200 12.500 54.300 ;
        RECT 15.800 54.200 16.100 55.800 ;
        RECT 19.000 55.600 19.400 59.900 ;
        RECT 21.100 57.200 21.500 59.900 ;
        RECT 20.600 56.800 21.500 57.200 ;
        RECT 21.800 56.800 22.200 57.200 ;
        RECT 21.100 56.200 21.500 56.800 ;
        RECT 21.900 56.200 22.200 56.800 ;
        RECT 21.100 55.900 21.600 56.200 ;
        RECT 21.900 55.900 22.600 56.200 ;
        RECT 17.300 55.300 19.400 55.600 ;
        RECT 17.300 55.200 17.700 55.300 ;
        RECT 18.100 54.900 18.500 55.000 ;
        RECT 16.600 54.600 18.500 54.900 ;
        RECT 16.600 54.500 17.000 54.600 ;
        RECT 10.600 53.900 16.100 54.200 ;
        RECT 10.600 53.800 11.400 53.900 ;
        RECT 7.900 53.300 9.800 53.600 ;
        RECT 7.900 53.200 8.300 53.300 ;
        RECT 2.200 52.100 2.600 52.500 ;
        RECT 3.000 52.400 3.400 53.200 ;
        RECT 3.900 52.700 4.300 52.800 ;
        RECT 3.900 52.400 5.300 52.700 ;
        RECT 5.000 52.100 5.300 52.400 ;
        RECT 7.000 52.100 7.400 52.500 ;
        RECT 2.200 51.800 3.200 52.100 ;
        RECT 2.800 51.100 3.200 51.800 ;
        RECT 5.000 51.100 5.400 52.100 ;
        RECT 7.000 51.800 7.700 52.100 ;
        RECT 7.100 51.100 7.700 51.800 ;
        RECT 9.400 51.100 9.800 53.300 ;
        RECT 10.200 51.100 10.600 53.500 ;
        RECT 12.700 52.800 13.000 53.900 ;
        RECT 15.500 53.800 15.900 53.900 ;
        RECT 19.000 53.600 19.400 55.300 ;
        RECT 19.800 55.100 20.200 55.200 ;
        RECT 20.600 55.100 21.000 55.200 ;
        RECT 19.800 54.800 21.000 55.100 ;
        RECT 20.600 54.400 21.000 54.800 ;
        RECT 21.300 54.200 21.600 55.900 ;
        RECT 22.200 55.800 22.600 55.900 ;
        RECT 23.000 55.800 23.400 56.600 ;
        RECT 22.200 55.100 22.500 55.800 ;
        RECT 23.800 55.100 24.200 59.900 ;
        RECT 25.400 55.700 25.800 59.900 ;
        RECT 27.600 58.200 28.000 59.900 ;
        RECT 27.000 57.900 28.000 58.200 ;
        RECT 29.800 57.900 30.200 59.900 ;
        RECT 31.900 57.900 32.500 59.900 ;
        RECT 27.000 57.500 27.400 57.900 ;
        RECT 29.800 57.600 30.100 57.900 ;
        RECT 28.700 57.300 30.500 57.600 ;
        RECT 31.800 57.500 32.200 57.900 ;
        RECT 28.700 57.200 29.100 57.300 ;
        RECT 30.100 57.200 30.500 57.300 ;
        RECT 34.200 57.100 34.600 59.900 ;
        RECT 35.000 57.100 35.400 57.200 ;
        RECT 27.000 56.500 27.400 56.600 ;
        RECT 29.300 56.500 29.700 56.600 ;
        RECT 27.000 56.200 29.700 56.500 ;
        RECT 30.000 56.500 31.100 56.800 ;
        RECT 30.000 55.900 30.300 56.500 ;
        RECT 30.700 56.400 31.100 56.500 ;
        RECT 31.900 56.600 32.600 57.000 ;
        RECT 34.200 56.800 35.400 57.100 ;
        RECT 31.900 56.100 32.200 56.600 ;
        RECT 27.900 55.700 30.300 55.900 ;
        RECT 25.400 55.600 30.300 55.700 ;
        RECT 31.000 55.800 32.200 56.100 ;
        RECT 25.400 55.500 28.300 55.600 ;
        RECT 25.400 55.400 28.200 55.500 ;
        RECT 28.600 55.100 29.000 55.200 ;
        RECT 29.400 55.100 29.800 55.200 ;
        RECT 22.200 54.800 24.200 55.100 ;
        RECT 19.800 54.100 20.200 54.200 ;
        RECT 19.800 53.800 20.600 54.100 ;
        RECT 21.300 53.800 22.600 54.200 ;
        RECT 20.200 53.600 20.600 53.800 ;
        RECT 17.500 53.300 19.400 53.600 ;
        RECT 17.500 53.200 17.900 53.300 ;
        RECT 11.800 52.100 12.200 52.500 ;
        RECT 12.600 52.400 13.000 52.800 ;
        RECT 13.500 52.700 13.900 52.800 ;
        RECT 13.500 52.400 14.900 52.700 ;
        RECT 14.600 52.100 14.900 52.400 ;
        RECT 16.600 52.100 17.000 52.500 ;
        RECT 11.800 51.800 12.800 52.100 ;
        RECT 12.400 51.100 12.800 51.800 ;
        RECT 14.600 51.100 15.000 52.100 ;
        RECT 16.600 51.800 17.300 52.100 ;
        RECT 16.700 51.100 17.300 51.800 ;
        RECT 19.000 51.100 19.400 53.300 ;
        RECT 19.900 53.100 21.700 53.300 ;
        RECT 22.200 53.100 22.500 53.800 ;
        RECT 23.800 53.100 24.200 54.800 ;
        RECT 26.500 54.800 29.800 55.100 ;
        RECT 26.500 54.700 26.900 54.800 ;
        RECT 27.300 54.200 27.700 54.300 ;
        RECT 31.000 54.200 31.300 55.800 ;
        RECT 34.200 55.600 34.600 56.800 ;
        RECT 32.500 55.300 34.600 55.600 ;
        RECT 32.500 55.200 32.900 55.300 ;
        RECT 33.300 54.900 33.700 55.000 ;
        RECT 31.800 54.600 33.700 54.900 ;
        RECT 31.800 54.500 32.200 54.600 ;
        RECT 24.600 53.400 25.000 54.200 ;
        RECT 25.800 53.900 31.300 54.200 ;
        RECT 34.200 54.100 34.600 55.300 ;
        RECT 35.800 55.100 36.200 59.900 ;
        RECT 37.800 56.800 38.200 57.200 ;
        RECT 36.600 55.800 37.000 56.600 ;
        RECT 37.800 56.200 38.100 56.800 ;
        RECT 38.500 56.200 38.900 59.900 ;
        RECT 41.900 59.200 42.300 59.900 ;
        RECT 41.400 58.800 42.300 59.200 ;
        RECT 37.400 55.900 38.100 56.200 ;
        RECT 38.400 55.900 38.900 56.200 ;
        RECT 41.900 56.200 42.300 58.800 ;
        RECT 42.600 56.800 43.000 57.200 ;
        RECT 42.700 56.200 43.000 56.800 ;
        RECT 41.900 55.900 42.400 56.200 ;
        RECT 42.700 55.900 43.400 56.200 ;
        RECT 37.400 55.800 37.800 55.900 ;
        RECT 37.400 55.100 37.700 55.800 ;
        RECT 38.400 55.200 38.700 55.900 ;
        RECT 35.800 54.800 37.700 55.100 ;
        RECT 38.200 54.800 38.700 55.200 ;
        RECT 35.000 54.100 35.400 54.200 ;
        RECT 25.800 53.800 26.600 53.900 ;
        RECT 19.800 53.000 21.800 53.100 ;
        RECT 19.800 51.100 20.200 53.000 ;
        RECT 21.400 51.100 21.800 53.000 ;
        RECT 22.200 51.100 22.600 53.100 ;
        RECT 23.300 52.800 24.200 53.100 ;
        RECT 23.300 51.100 23.700 52.800 ;
        RECT 25.400 51.100 25.800 53.500 ;
        RECT 27.900 53.200 28.200 53.900 ;
        RECT 30.700 53.800 31.100 53.900 ;
        RECT 34.200 53.800 35.400 54.100 ;
        RECT 34.200 53.600 34.600 53.800 ;
        RECT 32.700 53.300 34.600 53.600 ;
        RECT 35.000 53.400 35.400 53.800 ;
        RECT 32.700 53.200 33.100 53.300 ;
        RECT 27.000 52.100 27.400 52.500 ;
        RECT 27.800 52.400 28.200 53.200 ;
        RECT 28.700 52.700 29.100 52.800 ;
        RECT 28.700 52.400 30.100 52.700 ;
        RECT 29.800 52.100 30.100 52.400 ;
        RECT 31.800 52.100 32.200 52.500 ;
        RECT 27.000 51.800 28.000 52.100 ;
        RECT 27.600 51.100 28.000 51.800 ;
        RECT 29.800 51.100 30.200 52.100 ;
        RECT 31.800 51.800 32.500 52.100 ;
        RECT 31.900 51.100 32.500 51.800 ;
        RECT 34.200 51.100 34.600 53.300 ;
        RECT 35.800 53.100 36.200 54.800 ;
        RECT 38.400 54.200 38.700 54.800 ;
        RECT 39.000 54.400 39.400 55.200 ;
        RECT 41.400 54.400 41.800 55.200 ;
        RECT 42.100 54.200 42.400 55.900 ;
        RECT 43.000 55.800 43.400 55.900 ;
        RECT 43.800 55.700 44.200 59.900 ;
        RECT 46.000 58.200 46.400 59.900 ;
        RECT 45.400 57.900 46.400 58.200 ;
        RECT 48.200 57.900 48.600 59.900 ;
        RECT 50.300 57.900 50.900 59.900 ;
        RECT 45.400 57.500 45.800 57.900 ;
        RECT 48.200 57.600 48.500 57.900 ;
        RECT 47.100 57.300 48.900 57.600 ;
        RECT 50.200 57.500 50.600 57.900 ;
        RECT 47.100 57.200 47.500 57.300 ;
        RECT 48.500 57.200 48.900 57.300 ;
        RECT 45.400 56.500 45.800 56.600 ;
        RECT 47.700 56.500 48.100 56.600 ;
        RECT 45.400 56.200 48.100 56.500 ;
        RECT 48.400 56.500 49.500 56.800 ;
        RECT 48.400 55.900 48.700 56.500 ;
        RECT 49.100 56.400 49.500 56.500 ;
        RECT 50.300 56.600 51.000 57.000 ;
        RECT 50.300 56.100 50.600 56.600 ;
        RECT 46.300 55.700 48.700 55.900 ;
        RECT 43.800 55.600 48.700 55.700 ;
        RECT 49.400 55.800 50.600 56.100 ;
        RECT 43.800 55.500 46.700 55.600 ;
        RECT 43.800 55.400 46.600 55.500 ;
        RECT 47.000 55.100 47.400 55.200 ;
        RECT 44.900 54.800 47.400 55.100 ;
        RECT 44.900 54.700 45.300 54.800 ;
        RECT 45.700 54.200 46.100 54.300 ;
        RECT 49.400 54.200 49.700 55.800 ;
        RECT 52.600 55.600 53.000 59.900 ;
        RECT 56.300 57.200 56.700 59.900 ;
        RECT 55.800 56.800 56.700 57.200 ;
        RECT 57.000 56.800 57.400 57.200 ;
        RECT 56.300 56.200 56.700 56.800 ;
        RECT 57.100 56.200 57.400 56.800 ;
        RECT 56.300 55.900 56.800 56.200 ;
        RECT 57.100 55.900 57.800 56.200 ;
        RECT 50.900 55.300 53.000 55.600 ;
        RECT 50.900 55.200 51.300 55.300 ;
        RECT 51.700 54.900 52.100 55.000 ;
        RECT 50.200 54.600 52.100 54.900 ;
        RECT 50.200 54.500 50.600 54.600 ;
        RECT 37.400 53.800 38.700 54.200 ;
        RECT 39.800 54.100 40.200 54.200 ;
        RECT 39.400 53.800 40.200 54.100 ;
        RECT 40.600 54.100 41.000 54.200 ;
        RECT 40.600 53.800 41.400 54.100 ;
        RECT 42.100 53.800 43.400 54.200 ;
        RECT 44.200 53.900 49.700 54.200 ;
        RECT 44.200 53.800 45.000 53.900 ;
        RECT 46.200 53.800 46.600 53.900 ;
        RECT 49.100 53.800 49.500 53.900 ;
        RECT 37.500 53.100 37.800 53.800 ;
        RECT 39.400 53.600 39.800 53.800 ;
        RECT 41.000 53.600 41.400 53.800 ;
        RECT 38.300 53.100 40.100 53.300 ;
        RECT 40.700 53.100 42.500 53.300 ;
        RECT 43.000 53.100 43.300 53.800 ;
        RECT 35.800 52.800 36.700 53.100 ;
        RECT 36.300 51.100 36.700 52.800 ;
        RECT 37.400 51.100 37.800 53.100 ;
        RECT 38.200 53.000 40.200 53.100 ;
        RECT 38.200 51.100 38.600 53.000 ;
        RECT 39.800 51.100 40.200 53.000 ;
        RECT 40.600 53.000 42.600 53.100 ;
        RECT 40.600 51.100 41.000 53.000 ;
        RECT 42.200 51.100 42.600 53.000 ;
        RECT 43.000 51.100 43.400 53.100 ;
        RECT 43.800 51.100 44.200 53.500 ;
        RECT 46.300 52.800 46.600 53.800 ;
        RECT 52.600 53.600 53.000 55.300 ;
        RECT 55.800 54.400 56.200 55.200 ;
        RECT 56.500 54.200 56.800 55.900 ;
        RECT 57.400 55.800 57.800 55.900 ;
        RECT 58.200 55.800 58.600 56.600 ;
        RECT 57.400 55.100 57.700 55.800 ;
        RECT 59.000 55.100 59.400 59.900 ;
        RECT 61.700 59.200 62.100 59.900 ;
        RECT 61.700 58.800 62.600 59.200 ;
        RECT 61.000 56.800 61.400 57.200 ;
        RECT 61.000 56.200 61.300 56.800 ;
        RECT 61.700 56.200 62.100 58.800 ;
        RECT 60.600 55.900 61.300 56.200 ;
        RECT 61.600 55.900 62.100 56.200 ;
        RECT 63.800 56.200 64.200 59.900 ;
        RECT 65.400 56.200 65.800 59.900 ;
        RECT 63.800 55.900 65.800 56.200 ;
        RECT 66.200 55.900 66.600 59.900 ;
        RECT 60.600 55.800 61.000 55.900 ;
        RECT 57.400 54.800 59.400 55.100 ;
        RECT 53.400 54.100 53.800 54.200 ;
        RECT 55.000 54.100 55.400 54.200 ;
        RECT 53.400 53.800 55.800 54.100 ;
        RECT 56.500 53.800 57.800 54.200 ;
        RECT 55.400 53.600 55.800 53.800 ;
        RECT 51.100 53.300 53.000 53.600 ;
        RECT 51.100 53.200 51.500 53.300 ;
        RECT 45.400 52.100 45.800 52.500 ;
        RECT 46.200 52.400 46.600 52.800 ;
        RECT 47.100 52.700 47.500 52.800 ;
        RECT 47.100 52.400 48.500 52.700 ;
        RECT 48.200 52.100 48.500 52.400 ;
        RECT 50.200 52.100 50.600 52.500 ;
        RECT 45.400 51.800 46.400 52.100 ;
        RECT 46.000 51.100 46.400 51.800 ;
        RECT 48.200 51.100 48.600 52.100 ;
        RECT 50.200 51.800 50.900 52.100 ;
        RECT 50.300 51.100 50.900 51.800 ;
        RECT 52.600 51.100 53.000 53.300 ;
        RECT 55.100 53.100 56.900 53.300 ;
        RECT 57.400 53.100 57.700 53.800 ;
        RECT 59.000 53.100 59.400 54.800 ;
        RECT 61.600 54.200 61.900 55.900 ;
        RECT 64.200 55.200 64.600 55.400 ;
        RECT 66.200 55.200 66.500 55.900 ;
        RECT 67.000 55.700 67.400 59.900 ;
        RECT 69.200 58.200 69.600 59.900 ;
        RECT 68.600 57.900 69.600 58.200 ;
        RECT 71.400 57.900 71.800 59.900 ;
        RECT 73.500 57.900 74.100 59.900 ;
        RECT 68.600 57.500 69.000 57.900 ;
        RECT 71.400 57.600 71.700 57.900 ;
        RECT 70.300 57.300 72.100 57.600 ;
        RECT 73.400 57.500 73.800 57.900 ;
        RECT 70.300 57.200 70.700 57.300 ;
        RECT 71.700 57.200 72.100 57.300 ;
        RECT 68.600 56.500 69.000 56.600 ;
        RECT 70.900 56.500 71.300 56.600 ;
        RECT 68.600 56.200 71.300 56.500 ;
        RECT 71.600 56.500 72.700 56.800 ;
        RECT 71.600 55.900 71.900 56.500 ;
        RECT 72.300 56.400 72.700 56.500 ;
        RECT 73.500 56.600 74.200 57.000 ;
        RECT 73.500 56.100 73.800 56.600 ;
        RECT 69.500 55.700 71.900 55.900 ;
        RECT 67.000 55.600 71.900 55.700 ;
        RECT 72.600 55.800 73.800 56.100 ;
        RECT 67.000 55.500 69.900 55.600 ;
        RECT 67.000 55.400 69.800 55.500 ;
        RECT 62.200 54.400 62.600 55.200 ;
        RECT 63.000 55.100 63.400 55.200 ;
        RECT 63.800 55.100 64.600 55.200 ;
        RECT 63.000 54.900 64.600 55.100 ;
        RECT 65.400 54.900 66.600 55.200 ;
        RECT 70.200 55.100 70.600 55.200 ;
        RECT 63.000 54.800 64.200 54.900 ;
        RECT 65.400 54.800 65.800 54.900 ;
        RECT 66.200 54.800 66.600 54.900 ;
        RECT 68.100 54.800 70.600 55.100 ;
        RECT 59.800 53.400 60.200 54.200 ;
        RECT 60.600 53.800 61.900 54.200 ;
        RECT 63.000 54.100 63.400 54.200 ;
        RECT 62.600 53.800 63.400 54.100 ;
        RECT 64.600 53.800 65.000 54.600 ;
        RECT 60.700 53.100 61.000 53.800 ;
        RECT 62.600 53.600 63.000 53.800 ;
        RECT 61.500 53.100 63.300 53.300 ;
        RECT 65.400 53.100 65.700 54.800 ;
        RECT 68.100 54.700 68.500 54.800 ;
        RECT 68.900 54.200 69.300 54.300 ;
        RECT 72.600 54.200 72.900 55.800 ;
        RECT 75.800 55.600 76.200 59.900 ;
        RECT 77.900 56.200 78.300 59.900 ;
        RECT 78.600 56.800 79.000 57.200 ;
        RECT 78.700 56.200 79.000 56.800 ;
        RECT 77.400 55.800 78.400 56.200 ;
        RECT 78.700 55.900 79.400 56.200 ;
        RECT 74.100 55.300 76.200 55.600 ;
        RECT 74.100 55.200 74.500 55.300 ;
        RECT 74.900 54.900 75.300 55.000 ;
        RECT 73.400 54.600 75.300 54.900 ;
        RECT 73.400 54.500 73.800 54.600 ;
        RECT 67.400 53.900 72.900 54.200 ;
        RECT 67.400 53.800 68.200 53.900 ;
        RECT 55.000 53.000 57.000 53.100 ;
        RECT 55.000 51.100 55.400 53.000 ;
        RECT 56.600 51.100 57.000 53.000 ;
        RECT 57.400 51.100 57.800 53.100 ;
        RECT 58.500 52.800 59.400 53.100 ;
        RECT 58.500 51.100 58.900 52.800 ;
        RECT 60.600 51.100 61.000 53.100 ;
        RECT 61.400 53.000 63.400 53.100 ;
        RECT 61.400 51.100 61.800 53.000 ;
        RECT 63.000 51.100 63.400 53.000 ;
        RECT 65.400 51.100 65.800 53.100 ;
        RECT 66.200 52.800 66.600 53.200 ;
        RECT 66.100 52.400 66.500 52.800 ;
        RECT 67.000 51.100 67.400 53.500 ;
        RECT 69.500 52.800 69.800 53.900 ;
        RECT 71.000 53.800 71.400 53.900 ;
        RECT 72.300 53.800 72.700 53.900 ;
        RECT 75.800 53.600 76.200 55.300 ;
        RECT 77.400 54.400 77.800 55.200 ;
        RECT 78.100 54.200 78.400 55.800 ;
        RECT 79.000 55.800 79.400 55.900 ;
        RECT 79.800 55.800 80.200 56.600 ;
        RECT 79.000 55.100 79.300 55.800 ;
        RECT 80.600 55.100 81.000 59.900 ;
        RECT 82.200 55.900 82.600 59.900 ;
        RECT 83.000 56.200 83.400 59.900 ;
        RECT 84.600 56.200 85.000 59.900 ;
        RECT 86.500 59.200 86.900 59.900 ;
        RECT 86.500 58.800 87.400 59.200 ;
        RECT 85.800 56.800 86.200 57.200 ;
        RECT 85.800 56.200 86.100 56.800 ;
        RECT 86.500 56.200 86.900 58.800 ;
        RECT 83.000 55.900 85.000 56.200 ;
        RECT 85.400 55.900 86.100 56.200 ;
        RECT 86.400 55.900 86.900 56.200 ;
        RECT 89.900 56.200 90.300 59.900 ;
        RECT 90.600 56.800 91.000 57.200 ;
        RECT 90.700 56.200 91.000 56.800 ;
        RECT 89.900 55.900 90.400 56.200 ;
        RECT 90.700 55.900 91.400 56.200 ;
        RECT 82.300 55.200 82.600 55.900 ;
        RECT 85.400 55.800 85.800 55.900 ;
        RECT 84.200 55.200 84.600 55.400 ;
        RECT 79.000 54.800 81.000 55.100 ;
        RECT 82.200 54.900 83.400 55.200 ;
        RECT 84.200 54.900 85.000 55.200 ;
        RECT 82.200 54.800 82.600 54.900 ;
        RECT 76.600 54.100 77.000 54.200 ;
        RECT 76.600 53.800 77.400 54.100 ;
        RECT 78.100 53.800 79.400 54.200 ;
        RECT 77.000 53.600 77.400 53.800 ;
        RECT 74.300 53.300 76.200 53.600 ;
        RECT 74.300 53.200 74.700 53.300 ;
        RECT 68.600 52.100 69.000 52.500 ;
        RECT 69.400 52.400 69.800 52.800 ;
        RECT 70.300 52.700 70.700 52.800 ;
        RECT 70.300 52.400 71.700 52.700 ;
        RECT 71.400 52.100 71.700 52.400 ;
        RECT 73.400 52.100 73.800 52.500 ;
        RECT 68.600 51.800 69.600 52.100 ;
        RECT 69.200 51.100 69.600 51.800 ;
        RECT 71.400 51.100 71.800 52.100 ;
        RECT 73.400 51.800 74.100 52.100 ;
        RECT 73.500 51.100 74.100 51.800 ;
        RECT 75.800 51.100 76.200 53.300 ;
        RECT 76.700 53.100 78.500 53.300 ;
        RECT 79.000 53.100 79.300 53.800 ;
        RECT 80.600 53.100 81.000 54.800 ;
        RECT 81.400 53.400 81.800 54.200 ;
        RECT 83.100 53.200 83.400 54.900 ;
        RECT 84.600 54.800 85.000 54.900 ;
        RECT 83.800 53.800 84.200 54.600 ;
        RECT 86.400 54.200 86.700 55.900 ;
        RECT 87.000 54.400 87.400 55.200 ;
        RECT 89.400 54.400 89.800 55.200 ;
        RECT 90.100 54.200 90.400 55.900 ;
        RECT 91.000 55.800 91.400 55.900 ;
        RECT 91.800 55.800 92.200 56.600 ;
        RECT 91.000 55.100 91.300 55.800 ;
        RECT 92.600 55.100 93.000 59.900 ;
        RECT 94.200 55.700 94.600 59.900 ;
        RECT 96.400 58.200 96.800 59.900 ;
        RECT 95.800 57.900 96.800 58.200 ;
        RECT 98.600 57.900 99.000 59.900 ;
        RECT 100.700 57.900 101.300 59.900 ;
        RECT 95.800 57.500 96.200 57.900 ;
        RECT 98.600 57.600 98.900 57.900 ;
        RECT 97.500 57.300 99.300 57.600 ;
        RECT 100.600 57.500 101.000 57.900 ;
        RECT 97.500 57.200 97.900 57.300 ;
        RECT 98.900 57.200 99.300 57.300 ;
        RECT 95.800 56.500 96.200 56.600 ;
        RECT 98.100 56.500 98.500 56.600 ;
        RECT 95.800 56.200 98.500 56.500 ;
        RECT 98.800 56.500 99.900 56.800 ;
        RECT 98.800 55.900 99.100 56.500 ;
        RECT 99.500 56.400 99.900 56.500 ;
        RECT 100.700 56.600 101.400 57.000 ;
        RECT 100.700 56.100 101.000 56.600 ;
        RECT 96.700 55.700 99.100 55.900 ;
        RECT 94.200 55.600 99.100 55.700 ;
        RECT 99.800 55.800 101.000 56.100 ;
        RECT 94.200 55.500 97.100 55.600 ;
        RECT 94.200 55.400 97.000 55.500 ;
        RECT 99.800 55.200 100.100 55.800 ;
        RECT 103.000 55.600 103.400 59.900 ;
        RECT 106.500 59.200 106.900 59.900 ;
        RECT 106.500 58.800 107.400 59.200 ;
        RECT 105.800 56.800 106.200 57.200 ;
        RECT 105.800 56.200 106.100 56.800 ;
        RECT 106.500 56.200 106.900 58.800 ;
        RECT 104.600 56.100 105.000 56.200 ;
        RECT 105.400 56.100 106.100 56.200 ;
        RECT 104.600 55.900 106.100 56.100 ;
        RECT 106.400 55.900 106.900 56.200 ;
        RECT 104.600 55.800 105.800 55.900 ;
        RECT 101.300 55.300 103.400 55.600 ;
        RECT 101.300 55.200 101.700 55.300 ;
        RECT 97.400 55.100 97.800 55.200 ;
        RECT 91.000 54.800 93.000 55.100 ;
        RECT 85.400 53.800 86.700 54.200 ;
        RECT 87.800 54.100 88.200 54.200 ;
        RECT 87.400 53.800 88.200 54.100 ;
        RECT 88.600 54.100 89.000 54.200 ;
        RECT 90.100 54.100 91.400 54.200 ;
        RECT 91.800 54.100 92.200 54.200 ;
        RECT 88.600 53.800 89.400 54.100 ;
        RECT 90.100 53.800 92.200 54.100 ;
        RECT 76.600 53.000 78.600 53.100 ;
        RECT 76.600 51.100 77.000 53.000 ;
        RECT 78.200 51.100 78.600 53.000 ;
        RECT 79.000 51.100 79.400 53.100 ;
        RECT 80.100 52.800 81.000 53.100 ;
        RECT 82.200 52.800 82.600 53.200 ;
        RECT 80.100 51.100 80.500 52.800 ;
        RECT 82.300 52.400 82.700 52.800 ;
        RECT 83.000 51.100 83.400 53.200 ;
        RECT 85.500 53.100 85.800 53.800 ;
        RECT 87.400 53.600 87.800 53.800 ;
        RECT 89.000 53.600 89.400 53.800 ;
        RECT 86.300 53.100 88.100 53.300 ;
        RECT 88.700 53.100 90.500 53.300 ;
        RECT 91.000 53.100 91.300 53.800 ;
        RECT 92.600 53.100 93.000 54.800 ;
        RECT 95.300 54.800 97.800 55.100 ;
        RECT 99.800 54.800 100.200 55.200 ;
        RECT 102.100 54.900 102.500 55.000 ;
        RECT 95.300 54.700 95.700 54.800 ;
        RECT 96.600 54.700 97.000 54.800 ;
        RECT 96.100 54.200 96.500 54.300 ;
        RECT 99.800 54.200 100.100 54.800 ;
        RECT 100.600 54.600 102.500 54.900 ;
        RECT 100.600 54.500 101.000 54.600 ;
        RECT 93.400 53.400 93.800 54.200 ;
        RECT 94.600 53.900 100.100 54.200 ;
        RECT 94.600 53.800 95.400 53.900 ;
        RECT 85.400 51.100 85.800 53.100 ;
        RECT 86.200 53.000 88.200 53.100 ;
        RECT 86.200 51.100 86.600 53.000 ;
        RECT 87.800 51.100 88.200 53.000 ;
        RECT 88.600 53.000 90.600 53.100 ;
        RECT 88.600 51.100 89.000 53.000 ;
        RECT 90.200 51.100 90.600 53.000 ;
        RECT 91.000 51.100 91.400 53.100 ;
        RECT 92.100 52.800 93.000 53.100 ;
        RECT 92.100 51.100 92.500 52.800 ;
        RECT 94.200 51.100 94.600 53.500 ;
        RECT 96.700 52.800 97.000 53.900 ;
        RECT 99.500 53.800 99.900 53.900 ;
        RECT 103.000 53.600 103.400 55.300 ;
        RECT 106.400 54.200 106.700 55.900 ;
        RECT 107.000 55.100 107.400 55.200 ;
        RECT 108.600 55.100 109.000 59.900 ;
        RECT 107.000 54.800 109.000 55.100 ;
        RECT 107.000 54.400 107.400 54.800 ;
        RECT 105.400 53.800 106.700 54.200 ;
        RECT 107.800 54.100 108.200 54.200 ;
        RECT 107.400 53.800 108.200 54.100 ;
        RECT 101.500 53.300 103.400 53.600 ;
        RECT 101.500 53.200 101.900 53.300 ;
        RECT 95.800 52.100 96.200 52.500 ;
        RECT 96.600 52.400 97.000 52.800 ;
        RECT 97.500 52.700 97.900 52.800 ;
        RECT 97.500 52.400 98.900 52.700 ;
        RECT 98.600 52.100 98.900 52.400 ;
        RECT 100.600 52.100 101.000 52.500 ;
        RECT 95.800 51.800 96.800 52.100 ;
        RECT 96.400 51.100 96.800 51.800 ;
        RECT 98.600 51.100 99.000 52.100 ;
        RECT 100.600 51.800 101.300 52.100 ;
        RECT 100.700 51.100 101.300 51.800 ;
        RECT 103.000 51.100 103.400 53.300 ;
        RECT 105.500 53.100 105.800 53.800 ;
        RECT 107.400 53.600 107.800 53.800 ;
        RECT 106.300 53.100 108.100 53.300 ;
        RECT 105.400 51.100 105.800 53.100 ;
        RECT 106.200 53.000 108.200 53.100 ;
        RECT 106.200 51.100 106.600 53.000 ;
        RECT 107.800 51.100 108.200 53.000 ;
        RECT 108.600 51.100 109.000 54.800 ;
        RECT 111.000 55.100 111.400 59.900 ;
        RECT 113.000 56.800 113.400 57.200 ;
        RECT 111.800 55.800 112.200 56.600 ;
        RECT 113.000 56.200 113.300 56.800 ;
        RECT 113.700 56.200 114.100 59.900 ;
        RECT 112.600 55.900 113.300 56.200 ;
        RECT 113.600 55.900 114.100 56.200 ;
        RECT 115.800 56.200 116.200 59.900 ;
        RECT 117.400 56.200 117.800 59.900 ;
        RECT 115.800 55.900 117.800 56.200 ;
        RECT 118.200 55.900 118.600 59.900 ;
        RECT 112.600 55.800 113.000 55.900 ;
        RECT 112.600 55.100 112.900 55.800 ;
        RECT 111.000 54.800 112.900 55.100 ;
        RECT 110.200 54.100 110.600 54.200 ;
        RECT 109.400 53.800 110.600 54.100 ;
        RECT 109.400 53.200 109.700 53.800 ;
        RECT 110.200 53.400 110.600 53.800 ;
        RECT 109.400 52.400 109.800 53.200 ;
        RECT 111.000 53.100 111.400 54.800 ;
        RECT 113.600 54.200 113.900 55.900 ;
        RECT 116.200 55.200 116.600 55.400 ;
        RECT 118.200 55.200 118.500 55.900 ;
        RECT 119.000 55.600 119.400 59.900 ;
        RECT 121.100 57.900 121.700 59.900 ;
        RECT 123.400 57.900 123.800 59.900 ;
        RECT 125.600 58.200 126.000 59.900 ;
        RECT 125.600 57.900 126.600 58.200 ;
        RECT 121.400 57.500 121.800 57.900 ;
        RECT 123.500 57.600 123.800 57.900 ;
        RECT 123.100 57.300 124.900 57.600 ;
        RECT 126.200 57.500 126.600 57.900 ;
        RECT 123.100 57.200 123.500 57.300 ;
        RECT 124.500 57.200 124.900 57.300 ;
        RECT 121.000 56.600 121.700 57.000 ;
        RECT 121.400 56.100 121.700 56.600 ;
        RECT 122.500 56.500 123.600 56.800 ;
        RECT 122.500 56.400 122.900 56.500 ;
        RECT 121.400 55.800 122.600 56.100 ;
        RECT 119.000 55.300 121.100 55.600 ;
        RECT 114.200 54.400 114.600 55.200 ;
        RECT 115.800 54.900 116.600 55.200 ;
        RECT 117.400 54.900 118.600 55.200 ;
        RECT 115.800 54.800 116.200 54.900 ;
        RECT 112.600 53.800 113.900 54.200 ;
        RECT 115.000 54.100 115.400 54.200 ;
        RECT 114.600 53.800 115.400 54.100 ;
        RECT 116.600 53.800 117.000 54.600 ;
        RECT 112.700 53.100 113.000 53.800 ;
        RECT 114.600 53.600 115.000 53.800 ;
        RECT 113.500 53.100 115.300 53.300 ;
        RECT 117.400 53.100 117.700 54.900 ;
        RECT 118.200 54.800 118.600 54.900 ;
        RECT 119.000 53.600 119.400 55.300 ;
        RECT 120.700 55.200 121.100 55.300 ;
        RECT 119.900 54.900 120.300 55.000 ;
        RECT 119.900 54.600 121.800 54.900 ;
        RECT 121.400 54.500 121.800 54.600 ;
        RECT 122.300 54.200 122.600 55.800 ;
        RECT 123.300 55.900 123.600 56.500 ;
        RECT 123.900 56.500 124.300 56.600 ;
        RECT 126.200 56.500 126.600 56.600 ;
        RECT 123.900 56.200 126.600 56.500 ;
        RECT 123.300 55.700 125.700 55.900 ;
        RECT 127.800 55.700 128.200 59.900 ;
        RECT 129.900 56.200 130.300 59.900 ;
        RECT 130.600 56.800 131.000 57.200 ;
        RECT 130.700 56.200 131.000 56.800 ;
        RECT 129.900 55.900 130.400 56.200 ;
        RECT 130.700 55.900 131.400 56.200 ;
        RECT 123.300 55.600 128.200 55.700 ;
        RECT 125.300 55.500 128.200 55.600 ;
        RECT 125.400 55.400 128.200 55.500 ;
        RECT 130.100 55.200 130.400 55.900 ;
        RECT 131.000 55.800 131.400 55.900 ;
        RECT 131.800 55.800 132.200 56.600 ;
        RECT 123.800 55.100 124.200 55.200 ;
        RECT 124.600 55.100 125.000 55.200 ;
        RECT 123.800 54.800 127.100 55.100 ;
        RECT 126.700 54.700 127.100 54.800 ;
        RECT 129.400 54.400 129.800 55.200 ;
        RECT 130.100 54.800 130.600 55.200 ;
        RECT 131.000 55.100 131.300 55.800 ;
        RECT 132.600 55.100 133.000 59.900 ;
        RECT 134.200 55.700 134.600 59.900 ;
        RECT 136.400 58.200 136.800 59.900 ;
        RECT 135.800 57.900 136.800 58.200 ;
        RECT 138.600 57.900 139.000 59.900 ;
        RECT 140.700 57.900 141.300 59.900 ;
        RECT 135.800 57.500 136.200 57.900 ;
        RECT 138.600 57.600 138.900 57.900 ;
        RECT 137.500 57.300 139.300 57.600 ;
        RECT 140.600 57.500 141.000 57.900 ;
        RECT 137.500 57.200 137.900 57.300 ;
        RECT 138.900 57.200 139.300 57.300 ;
        RECT 135.800 56.500 136.200 56.600 ;
        RECT 138.100 56.500 138.500 56.600 ;
        RECT 135.800 56.200 138.500 56.500 ;
        RECT 138.800 56.500 139.900 56.800 ;
        RECT 138.800 55.900 139.100 56.500 ;
        RECT 139.500 56.400 139.900 56.500 ;
        RECT 140.700 56.600 141.400 57.000 ;
        RECT 140.700 56.100 141.000 56.600 ;
        RECT 136.700 55.700 139.100 55.900 ;
        RECT 134.200 55.600 139.100 55.700 ;
        RECT 139.800 55.800 141.000 56.100 ;
        RECT 134.200 55.500 137.100 55.600 ;
        RECT 134.200 55.400 137.000 55.500 ;
        RECT 139.800 55.200 140.100 55.800 ;
        RECT 143.000 55.600 143.400 59.900 ;
        RECT 143.800 56.200 144.200 59.900 ;
        RECT 145.400 56.400 145.800 59.900 ;
        RECT 143.800 55.900 145.100 56.200 ;
        RECT 145.400 55.900 145.900 56.400 ;
        RECT 141.300 55.300 143.400 55.600 ;
        RECT 141.300 55.200 141.700 55.300 ;
        RECT 137.400 55.100 137.800 55.200 ;
        RECT 131.000 54.800 133.000 55.100 ;
        RECT 125.900 54.200 126.300 54.300 ;
        RECT 130.100 54.200 130.400 54.800 ;
        RECT 122.300 53.900 127.800 54.200 ;
        RECT 122.500 53.800 122.900 53.900 ;
        RECT 124.600 53.800 125.000 53.900 ;
        RECT 119.000 53.300 120.900 53.600 ;
        RECT 111.000 52.800 111.900 53.100 ;
        RECT 111.500 51.100 111.900 52.800 ;
        RECT 112.600 51.100 113.000 53.100 ;
        RECT 113.400 53.000 115.400 53.100 ;
        RECT 113.400 51.100 113.800 53.000 ;
        RECT 115.000 51.100 115.400 53.000 ;
        RECT 117.400 51.100 117.800 53.100 ;
        RECT 118.200 52.800 118.600 53.200 ;
        RECT 118.100 52.400 118.500 52.800 ;
        RECT 119.000 51.100 119.400 53.300 ;
        RECT 120.500 53.200 120.900 53.300 ;
        RECT 125.400 52.800 125.700 53.900 ;
        RECT 127.000 53.800 127.800 53.900 ;
        RECT 128.600 54.100 129.000 54.200 ;
        RECT 128.600 53.800 129.400 54.100 ;
        RECT 130.100 53.800 131.400 54.200 ;
        RECT 129.000 53.600 129.400 53.800 ;
        RECT 124.500 52.700 124.900 52.800 ;
        RECT 121.400 52.100 121.800 52.500 ;
        RECT 123.500 52.400 124.900 52.700 ;
        RECT 125.400 52.400 125.800 52.800 ;
        RECT 123.500 52.100 123.800 52.400 ;
        RECT 126.200 52.100 126.600 52.500 ;
        RECT 121.100 51.800 121.800 52.100 ;
        RECT 121.100 51.100 121.700 51.800 ;
        RECT 123.400 51.100 123.800 52.100 ;
        RECT 125.600 51.800 126.600 52.100 ;
        RECT 125.600 51.100 126.000 51.800 ;
        RECT 127.800 51.100 128.200 53.500 ;
        RECT 128.700 53.100 130.500 53.300 ;
        RECT 131.000 53.100 131.300 53.800 ;
        RECT 132.600 53.100 133.000 54.800 ;
        RECT 135.300 54.800 137.800 55.100 ;
        RECT 139.800 54.800 140.200 55.200 ;
        RECT 142.100 54.900 142.500 55.000 ;
        RECT 135.300 54.700 135.700 54.800 ;
        RECT 136.600 54.700 137.000 54.800 ;
        RECT 136.100 54.200 136.500 54.300 ;
        RECT 139.800 54.200 140.100 54.800 ;
        RECT 140.600 54.600 142.500 54.900 ;
        RECT 140.600 54.500 141.000 54.600 ;
        RECT 133.400 53.400 133.800 54.200 ;
        RECT 134.600 53.900 140.100 54.200 ;
        RECT 134.600 53.800 135.400 53.900 ;
        RECT 128.600 53.000 130.600 53.100 ;
        RECT 128.600 51.100 129.000 53.000 ;
        RECT 130.200 51.100 130.600 53.000 ;
        RECT 131.000 51.100 131.400 53.100 ;
        RECT 132.100 52.800 133.000 53.100 ;
        RECT 132.100 51.100 132.500 52.800 ;
        RECT 134.200 51.100 134.600 53.500 ;
        RECT 136.700 52.800 137.000 53.900 ;
        RECT 139.500 53.800 139.900 53.900 ;
        RECT 141.400 53.600 141.800 54.200 ;
        RECT 143.000 53.600 143.400 55.300 ;
        RECT 143.800 54.800 144.300 55.200 ;
        RECT 143.900 54.400 144.300 54.800 ;
        RECT 144.800 54.900 145.100 55.900 ;
        RECT 144.800 54.500 145.300 54.900 ;
        RECT 144.800 53.700 145.100 54.500 ;
        RECT 145.600 54.200 145.900 55.900 ;
        RECT 145.400 53.800 145.900 54.200 ;
        RECT 141.400 53.300 143.400 53.600 ;
        RECT 141.500 53.200 141.900 53.300 ;
        RECT 135.800 52.100 136.200 52.500 ;
        RECT 136.600 52.400 137.000 52.800 ;
        RECT 137.500 52.700 137.900 52.800 ;
        RECT 137.500 52.400 138.900 52.700 ;
        RECT 138.600 52.100 138.900 52.400 ;
        RECT 140.600 52.100 141.000 52.500 ;
        RECT 135.800 51.800 136.800 52.100 ;
        RECT 136.400 51.100 136.800 51.800 ;
        RECT 138.600 51.100 139.000 52.100 ;
        RECT 140.600 51.800 141.300 52.100 ;
        RECT 140.700 51.100 141.300 51.800 ;
        RECT 143.000 51.100 143.400 53.300 ;
        RECT 143.800 53.400 145.100 53.700 ;
        RECT 143.800 51.100 144.200 53.400 ;
        RECT 145.600 53.100 145.900 53.800 ;
        RECT 145.400 52.800 145.900 53.100 ;
        RECT 147.000 55.600 147.400 59.900 ;
        RECT 149.100 57.900 149.700 59.900 ;
        RECT 151.400 57.900 151.800 59.900 ;
        RECT 153.600 58.200 154.000 59.900 ;
        RECT 153.600 57.900 154.600 58.200 ;
        RECT 149.400 57.500 149.800 57.900 ;
        RECT 151.500 57.600 151.800 57.900 ;
        RECT 151.100 57.300 152.900 57.600 ;
        RECT 154.200 57.500 154.600 57.900 ;
        RECT 151.100 57.200 151.500 57.300 ;
        RECT 152.500 57.200 152.900 57.300 ;
        RECT 149.000 56.600 149.700 57.000 ;
        RECT 149.400 56.100 149.700 56.600 ;
        RECT 150.500 56.500 151.600 56.800 ;
        RECT 150.500 56.400 150.900 56.500 ;
        RECT 149.400 55.800 150.600 56.100 ;
        RECT 147.000 55.300 149.100 55.600 ;
        RECT 147.000 53.600 147.400 55.300 ;
        RECT 148.700 55.200 149.100 55.300 ;
        RECT 150.300 55.200 150.600 55.800 ;
        RECT 151.300 55.900 151.600 56.500 ;
        RECT 151.900 56.500 152.300 56.600 ;
        RECT 154.200 56.500 154.600 56.600 ;
        RECT 151.900 56.200 154.600 56.500 ;
        RECT 151.300 55.700 153.700 55.900 ;
        RECT 155.800 55.700 156.200 59.900 ;
        RECT 151.300 55.600 156.200 55.700 ;
        RECT 153.300 55.500 156.200 55.600 ;
        RECT 153.400 55.400 156.200 55.500 ;
        RECT 147.900 54.900 148.300 55.000 ;
        RECT 147.900 54.600 149.800 54.900 ;
        RECT 150.200 54.800 150.600 55.200 ;
        RECT 152.600 55.100 153.000 55.200 ;
        RECT 158.200 55.100 158.600 59.900 ;
        RECT 159.000 55.800 159.400 56.200 ;
        RECT 159.000 55.100 159.300 55.800 ;
        RECT 152.600 54.800 155.100 55.100 ;
        RECT 149.400 54.500 149.800 54.600 ;
        RECT 150.300 54.200 150.600 54.800 ;
        RECT 153.400 54.700 153.800 54.800 ;
        RECT 154.700 54.700 155.100 54.800 ;
        RECT 158.200 54.800 159.300 55.100 ;
        RECT 159.800 55.600 160.200 59.900 ;
        RECT 161.900 57.900 162.500 59.900 ;
        RECT 164.200 57.900 164.600 59.900 ;
        RECT 166.400 58.200 166.800 59.900 ;
        RECT 166.400 57.900 167.400 58.200 ;
        RECT 162.200 57.500 162.600 57.900 ;
        RECT 164.300 57.600 164.600 57.900 ;
        RECT 163.900 57.300 165.700 57.600 ;
        RECT 167.000 57.500 167.400 57.900 ;
        RECT 163.900 57.200 164.300 57.300 ;
        RECT 165.300 57.200 165.700 57.300 ;
        RECT 161.800 56.600 162.500 57.000 ;
        RECT 162.200 56.100 162.500 56.600 ;
        RECT 163.300 56.500 164.400 56.800 ;
        RECT 163.300 56.400 163.700 56.500 ;
        RECT 162.200 55.800 163.400 56.100 ;
        RECT 159.800 55.300 161.900 55.600 ;
        RECT 153.900 54.200 154.300 54.300 ;
        RECT 150.300 54.100 155.800 54.200 ;
        RECT 156.600 54.100 157.000 54.200 ;
        RECT 150.300 53.900 157.000 54.100 ;
        RECT 150.500 53.800 150.900 53.900 ;
        RECT 147.000 53.300 148.900 53.600 ;
        RECT 145.400 51.100 145.800 52.800 ;
        RECT 147.000 51.100 147.400 53.300 ;
        RECT 148.500 53.200 148.900 53.300 ;
        RECT 153.400 52.800 153.700 53.900 ;
        RECT 155.000 53.800 157.000 53.900 ;
        RECT 152.500 52.700 152.900 52.800 ;
        RECT 149.400 52.100 149.800 52.500 ;
        RECT 151.500 52.400 152.900 52.700 ;
        RECT 153.400 52.400 153.800 52.800 ;
        RECT 151.500 52.100 151.800 52.400 ;
        RECT 154.200 52.100 154.600 52.500 ;
        RECT 149.100 51.800 149.800 52.100 ;
        RECT 149.100 51.100 149.700 51.800 ;
        RECT 151.400 51.100 151.800 52.100 ;
        RECT 153.600 51.800 154.600 52.100 ;
        RECT 153.600 51.100 154.000 51.800 ;
        RECT 155.800 51.100 156.200 53.500 ;
        RECT 158.200 51.100 158.600 54.800 ;
        RECT 159.800 53.600 160.200 55.300 ;
        RECT 161.500 55.200 161.900 55.300 ;
        RECT 160.700 54.900 161.100 55.000 ;
        RECT 160.700 54.600 162.600 54.900 ;
        RECT 162.200 54.500 162.600 54.600 ;
        RECT 163.100 54.200 163.400 55.800 ;
        RECT 164.100 55.900 164.400 56.500 ;
        RECT 164.700 56.500 165.100 56.600 ;
        RECT 167.000 56.500 167.400 56.600 ;
        RECT 164.700 56.200 167.400 56.500 ;
        RECT 164.100 55.700 166.500 55.900 ;
        RECT 168.600 55.700 169.000 59.900 ;
        RECT 164.100 55.600 169.000 55.700 ;
        RECT 166.100 55.500 169.000 55.600 ;
        RECT 169.400 57.500 169.800 59.500 ;
        RECT 169.400 55.800 169.700 57.500 ;
        RECT 171.500 56.400 171.900 59.900 ;
        RECT 171.500 56.100 172.300 56.400 ;
        RECT 169.400 55.500 171.300 55.800 ;
        RECT 166.200 55.400 169.000 55.500 ;
        RECT 165.400 55.100 165.800 55.200 ;
        RECT 165.400 54.800 167.900 55.100 ;
        RECT 166.200 54.700 166.600 54.800 ;
        RECT 167.500 54.700 167.900 54.800 ;
        RECT 169.400 54.400 169.800 55.200 ;
        RECT 170.200 54.400 170.600 55.200 ;
        RECT 171.000 54.500 171.300 55.500 ;
        RECT 166.700 54.200 167.100 54.300 ;
        RECT 163.100 53.900 168.600 54.200 ;
        RECT 171.000 54.100 171.700 54.500 ;
        RECT 172.000 54.200 172.300 56.100 ;
        RECT 174.200 56.200 174.600 59.900 ;
        RECT 175.800 56.200 176.200 59.900 ;
        RECT 174.200 55.900 176.200 56.200 ;
        RECT 176.600 55.900 177.000 59.900 ;
        RECT 177.800 56.800 178.200 57.200 ;
        RECT 177.800 56.200 178.100 56.800 ;
        RECT 178.500 56.200 178.900 59.900 ;
        RECT 177.400 55.900 178.100 56.200 ;
        RECT 178.400 55.900 178.900 56.200 ;
        RECT 172.600 55.100 173.000 55.600 ;
        RECT 174.600 55.200 175.000 55.400 ;
        RECT 176.600 55.200 176.900 55.900 ;
        RECT 177.400 55.800 177.800 55.900 ;
        RECT 173.400 55.100 173.800 55.200 ;
        RECT 172.600 54.800 173.800 55.100 ;
        RECT 174.200 54.900 175.000 55.200 ;
        RECT 175.800 54.900 177.000 55.200 ;
        RECT 174.200 54.800 174.600 54.900 ;
        RECT 171.000 53.900 171.500 54.100 ;
        RECT 163.300 53.800 163.700 53.900 ;
        RECT 165.400 53.800 165.800 53.900 ;
        RECT 159.800 53.300 161.700 53.600 ;
        RECT 159.000 53.100 159.400 53.200 ;
        RECT 159.800 53.100 160.200 53.300 ;
        RECT 161.300 53.200 161.700 53.300 ;
        RECT 159.000 52.800 160.200 53.100 ;
        RECT 166.200 52.800 166.500 53.900 ;
        RECT 167.800 53.800 168.600 53.900 ;
        RECT 169.400 53.600 171.500 53.900 ;
        RECT 172.000 53.800 173.000 54.200 ;
        RECT 175.000 53.800 175.400 54.600 ;
        RECT 159.000 52.400 159.400 52.800 ;
        RECT 159.800 51.100 160.200 52.800 ;
        RECT 165.300 52.700 165.700 52.800 ;
        RECT 162.200 52.100 162.600 52.500 ;
        RECT 164.300 52.400 165.700 52.700 ;
        RECT 166.200 52.400 166.600 52.800 ;
        RECT 164.300 52.100 164.600 52.400 ;
        RECT 167.000 52.100 167.400 52.500 ;
        RECT 161.900 51.800 162.600 52.100 ;
        RECT 161.900 51.100 162.500 51.800 ;
        RECT 164.200 51.100 164.600 52.100 ;
        RECT 166.400 51.800 167.400 52.100 ;
        RECT 166.400 51.100 166.800 51.800 ;
        RECT 168.600 51.100 169.000 53.500 ;
        RECT 169.400 52.500 169.700 53.600 ;
        RECT 172.000 53.500 172.300 53.800 ;
        RECT 171.900 53.300 172.300 53.500 ;
        RECT 171.500 53.000 172.300 53.300 ;
        RECT 175.800 53.100 176.100 54.900 ;
        RECT 176.600 54.800 177.000 54.900 ;
        RECT 178.400 54.200 178.700 55.900 ;
        RECT 180.600 55.700 181.000 59.900 ;
        RECT 182.800 58.200 183.200 59.900 ;
        RECT 182.200 57.900 183.200 58.200 ;
        RECT 185.000 57.900 185.400 59.900 ;
        RECT 187.100 57.900 187.700 59.900 ;
        RECT 182.200 57.500 182.600 57.900 ;
        RECT 185.000 57.600 185.300 57.900 ;
        RECT 183.900 57.300 185.700 57.600 ;
        RECT 187.000 57.500 187.400 57.900 ;
        RECT 183.900 57.200 184.300 57.300 ;
        RECT 185.300 57.200 185.700 57.300 ;
        RECT 182.200 56.500 182.600 56.600 ;
        RECT 184.500 56.500 184.900 56.600 ;
        RECT 182.200 56.200 184.900 56.500 ;
        RECT 185.200 56.500 186.300 56.800 ;
        RECT 185.200 55.900 185.500 56.500 ;
        RECT 185.900 56.400 186.300 56.500 ;
        RECT 187.100 56.600 187.800 57.000 ;
        RECT 187.100 56.100 187.400 56.600 ;
        RECT 183.100 55.700 185.500 55.900 ;
        RECT 180.600 55.600 185.500 55.700 ;
        RECT 186.200 55.800 187.400 56.100 ;
        RECT 180.600 55.500 183.500 55.600 ;
        RECT 180.600 55.400 183.400 55.500 ;
        RECT 179.000 54.400 179.400 55.200 ;
        RECT 183.800 55.100 184.200 55.200 ;
        RECT 181.700 54.800 184.200 55.100 ;
        RECT 181.700 54.700 182.100 54.800 ;
        RECT 183.000 54.700 183.400 54.800 ;
        RECT 182.500 54.200 182.900 54.300 ;
        RECT 186.200 54.200 186.500 55.800 ;
        RECT 189.400 55.600 189.800 59.900 ;
        RECT 187.700 55.300 189.800 55.600 ;
        RECT 187.700 55.200 188.100 55.300 ;
        RECT 188.500 54.900 188.900 55.000 ;
        RECT 187.000 54.600 188.900 54.900 ;
        RECT 187.000 54.500 187.400 54.600 ;
        RECT 177.400 53.800 178.700 54.200 ;
        RECT 179.800 54.100 180.200 54.200 ;
        RECT 179.400 53.800 180.200 54.100 ;
        RECT 181.000 53.900 186.500 54.200 ;
        RECT 181.000 53.800 181.800 53.900 ;
        RECT 176.600 53.100 177.000 53.200 ;
        RECT 177.500 53.100 177.800 53.800 ;
        RECT 179.400 53.600 179.800 53.800 ;
        RECT 178.300 53.100 180.100 53.300 ;
        RECT 171.500 52.800 172.200 53.000 ;
        RECT 169.400 51.500 169.800 52.500 ;
        RECT 171.500 51.500 171.900 52.800 ;
        RECT 175.800 51.100 176.200 53.100 ;
        RECT 176.600 52.800 177.800 53.100 ;
        RECT 176.500 52.400 176.900 52.800 ;
        RECT 177.400 51.100 177.800 52.800 ;
        RECT 178.200 53.000 180.200 53.100 ;
        RECT 178.200 51.100 178.600 53.000 ;
        RECT 179.800 51.100 180.200 53.000 ;
        RECT 180.600 51.100 181.000 53.500 ;
        RECT 183.100 52.800 183.400 53.900 ;
        RECT 185.900 53.800 186.300 53.900 ;
        RECT 189.400 53.600 189.800 55.300 ;
        RECT 187.900 53.300 189.800 53.600 ;
        RECT 187.900 53.200 188.300 53.300 ;
        RECT 189.400 53.100 189.800 53.300 ;
        RECT 190.200 53.100 190.600 53.200 ;
        RECT 189.400 52.800 190.600 53.100 ;
        RECT 182.200 52.100 182.600 52.500 ;
        RECT 183.000 52.400 183.400 52.800 ;
        RECT 183.900 52.700 184.300 52.800 ;
        RECT 183.900 52.400 185.300 52.700 ;
        RECT 185.000 52.100 185.300 52.400 ;
        RECT 187.000 52.100 187.400 52.500 ;
        RECT 182.200 51.800 183.200 52.100 ;
        RECT 182.800 51.100 183.200 51.800 ;
        RECT 185.000 51.100 185.400 52.100 ;
        RECT 187.000 51.800 187.700 52.100 ;
        RECT 187.100 51.100 187.700 51.800 ;
        RECT 189.400 51.100 189.800 52.800 ;
        RECT 190.200 52.400 190.600 52.800 ;
        RECT 191.000 51.100 191.400 59.900 ;
        RECT 191.800 55.800 192.200 56.600 ;
        RECT 192.600 53.100 193.000 59.900 ;
        RECT 194.200 56.200 194.600 59.900 ;
        RECT 195.800 56.200 196.200 59.900 ;
        RECT 194.200 55.900 196.200 56.200 ;
        RECT 196.600 55.900 197.000 59.900 ;
        RECT 197.700 56.300 198.100 59.900 ;
        RECT 197.700 55.900 198.600 56.300 ;
        RECT 194.600 55.200 195.000 55.400 ;
        RECT 196.600 55.200 196.900 55.900 ;
        RECT 193.400 55.100 193.800 55.200 ;
        RECT 194.200 55.100 195.000 55.200 ;
        RECT 193.400 54.900 195.000 55.100 ;
        RECT 195.800 54.900 197.000 55.200 ;
        RECT 193.400 54.800 194.600 54.900 ;
        RECT 194.200 54.100 194.600 54.200 ;
        RECT 195.000 54.100 195.400 54.600 ;
        RECT 194.200 53.800 195.400 54.100 ;
        RECT 192.100 52.800 193.000 53.100 ;
        RECT 195.800 53.100 196.100 54.900 ;
        RECT 196.600 54.800 197.000 54.900 ;
        RECT 197.400 54.800 197.800 55.600 ;
        RECT 198.200 54.200 198.500 55.900 ;
        RECT 199.800 55.800 200.200 56.600 ;
        RECT 199.000 55.100 199.400 55.200 ;
        RECT 200.600 55.100 201.000 59.900 ;
        RECT 202.200 55.900 202.600 59.900 ;
        RECT 203.000 56.200 203.400 59.900 ;
        RECT 204.600 56.200 205.000 59.900 ;
        RECT 203.000 55.900 205.000 56.200 ;
        RECT 202.300 55.200 202.600 55.900 ;
        RECT 204.200 55.200 204.600 55.400 ;
        RECT 199.000 54.800 201.000 55.100 ;
        RECT 202.200 54.900 203.400 55.200 ;
        RECT 204.200 54.900 205.000 55.200 ;
        RECT 202.200 54.800 202.600 54.900 ;
        RECT 198.200 53.800 198.600 54.200 ;
        RECT 196.600 53.100 197.000 53.200 ;
        RECT 198.200 53.100 198.500 53.800 ;
        RECT 192.100 51.100 192.500 52.800 ;
        RECT 195.800 51.100 196.200 53.100 ;
        RECT 196.600 52.800 198.500 53.100 ;
        RECT 196.500 52.400 196.900 52.800 ;
        RECT 198.200 52.100 198.500 52.800 ;
        RECT 199.000 52.400 199.400 53.200 ;
        RECT 200.600 53.100 201.000 54.800 ;
        RECT 200.100 52.800 201.000 53.100 ;
        RECT 202.200 52.800 202.600 53.200 ;
        RECT 203.100 53.100 203.400 54.900 ;
        RECT 204.600 54.800 205.000 54.900 ;
        RECT 203.800 53.800 204.200 54.600 ;
        RECT 198.200 51.100 198.600 52.100 ;
        RECT 200.100 51.100 200.500 52.800 ;
        RECT 202.300 52.400 202.700 52.800 ;
        RECT 203.000 51.100 203.400 53.100 ;
        RECT 1.400 47.600 1.800 49.900 ;
        RECT 3.000 47.600 3.400 49.900 ;
        RECT 4.600 47.600 5.000 49.900 ;
        RECT 6.200 47.600 6.600 49.900 ;
        RECT 8.600 48.900 9.000 49.900 ;
        RECT 7.800 47.800 8.200 48.600 ;
        RECT 8.700 48.100 9.000 48.900 ;
        RECT 10.300 48.200 10.700 48.600 ;
        RECT 10.200 48.100 10.600 48.200 ;
        RECT 8.600 47.800 10.600 48.100 ;
        RECT 11.000 47.900 11.400 49.900 ;
        RECT 14.700 48.200 15.100 49.900 ;
        RECT 1.400 47.200 2.300 47.600 ;
        RECT 3.000 47.200 4.100 47.600 ;
        RECT 4.600 47.200 5.700 47.600 ;
        RECT 6.200 47.200 7.400 47.600 ;
        RECT 8.700 47.200 9.000 47.800 ;
        RECT 1.900 46.900 2.300 47.200 ;
        RECT 3.700 46.900 4.100 47.200 ;
        RECT 5.300 46.900 5.700 47.200 ;
        RECT 1.900 46.500 3.200 46.900 ;
        RECT 3.700 46.500 4.900 46.900 ;
        RECT 5.300 46.500 6.600 46.900 ;
        RECT 1.900 45.800 2.300 46.500 ;
        RECT 3.700 45.800 4.100 46.500 ;
        RECT 5.300 45.800 5.700 46.500 ;
        RECT 7.000 45.800 7.400 47.200 ;
        RECT 8.600 46.800 9.000 47.200 ;
        RECT 1.400 45.400 2.300 45.800 ;
        RECT 3.000 45.400 4.100 45.800 ;
        RECT 4.600 45.400 5.700 45.800 ;
        RECT 6.200 45.400 7.400 45.800 ;
        RECT 1.400 41.100 1.800 45.400 ;
        RECT 3.000 41.100 3.400 45.400 ;
        RECT 4.600 41.100 5.000 45.400 ;
        RECT 6.200 41.100 6.600 45.400 ;
        RECT 8.700 45.100 9.000 46.800 ;
        RECT 9.400 45.400 9.800 46.200 ;
        RECT 10.200 46.100 10.600 46.200 ;
        RECT 11.100 46.100 11.400 47.900 ;
        RECT 14.200 47.900 15.100 48.200 ;
        RECT 15.800 47.900 16.200 49.900 ;
        RECT 16.600 48.000 17.000 49.900 ;
        RECT 18.200 48.000 18.600 49.900 ;
        RECT 16.600 47.900 18.600 48.000 ;
        RECT 19.000 48.000 19.400 49.900 ;
        RECT 20.600 48.000 21.000 49.900 ;
        RECT 19.000 47.900 21.000 48.000 ;
        RECT 21.400 47.900 21.800 49.900 ;
        RECT 22.500 48.200 22.900 49.900 ;
        RECT 22.500 47.900 23.400 48.200 ;
        RECT 11.800 47.100 12.200 47.200 ;
        RECT 12.600 47.100 13.000 47.200 ;
        RECT 11.800 46.800 13.000 47.100 ;
        RECT 13.400 46.800 13.800 47.600 ;
        RECT 11.800 46.400 12.200 46.800 ;
        RECT 12.600 46.100 13.000 46.200 ;
        RECT 10.200 45.800 11.400 46.100 ;
        RECT 12.200 45.800 13.000 46.100 ;
        RECT 14.200 46.100 14.600 47.900 ;
        RECT 15.900 47.200 16.200 47.900 ;
        RECT 16.700 47.700 18.500 47.900 ;
        RECT 19.100 47.700 20.900 47.900 ;
        RECT 17.800 47.200 18.200 47.400 ;
        RECT 19.400 47.200 19.800 47.400 ;
        RECT 21.400 47.200 21.700 47.900 ;
        RECT 15.800 46.800 17.100 47.200 ;
        RECT 17.800 47.100 18.600 47.200 ;
        RECT 19.000 47.100 19.800 47.200 ;
        RECT 17.800 46.900 19.800 47.100 ;
        RECT 20.500 47.100 21.800 47.200 ;
        RECT 22.200 47.100 22.600 47.200 ;
        RECT 18.200 46.800 19.400 46.900 ;
        RECT 20.500 46.800 22.600 47.100 ;
        RECT 14.200 45.800 16.100 46.100 ;
        RECT 10.300 45.100 10.600 45.800 ;
        RECT 12.200 45.600 12.600 45.800 ;
        RECT 8.600 44.700 9.500 45.100 ;
        RECT 9.100 41.100 9.500 44.700 ;
        RECT 10.200 41.100 10.600 45.100 ;
        RECT 11.000 44.800 13.000 45.100 ;
        RECT 11.000 41.100 11.400 44.800 ;
        RECT 12.600 41.100 13.000 44.800 ;
        RECT 14.200 41.100 14.600 45.800 ;
        RECT 15.800 45.200 16.100 45.800 ;
        RECT 15.000 44.400 15.400 45.200 ;
        RECT 15.800 45.100 16.200 45.200 ;
        RECT 16.800 45.100 17.100 46.800 ;
        RECT 17.400 45.800 17.800 46.600 ;
        RECT 18.200 46.100 18.600 46.200 ;
        RECT 19.800 46.100 20.200 46.600 ;
        RECT 18.200 45.800 20.200 46.100 ;
        RECT 20.500 45.100 20.800 46.800 ;
        RECT 23.000 46.100 23.400 47.900 ;
        RECT 23.800 46.800 24.200 47.600 ;
        RECT 24.600 47.500 25.000 49.900 ;
        RECT 26.800 49.200 27.200 49.900 ;
        RECT 26.200 48.900 27.200 49.200 ;
        RECT 29.000 48.900 29.400 49.900 ;
        RECT 31.100 49.200 31.700 49.900 ;
        RECT 31.000 48.900 31.700 49.200 ;
        RECT 26.200 48.500 26.600 48.900 ;
        RECT 29.000 48.600 29.300 48.900 ;
        RECT 27.000 48.200 27.400 48.600 ;
        RECT 27.900 48.300 29.300 48.600 ;
        RECT 31.000 48.500 31.400 48.900 ;
        RECT 27.900 48.200 28.300 48.300 ;
        RECT 25.000 47.100 25.800 47.200 ;
        RECT 27.100 47.100 27.400 48.200 ;
        RECT 31.900 47.700 32.300 47.800 ;
        RECT 33.400 47.700 33.800 49.900 ;
        RECT 34.200 48.000 34.600 49.900 ;
        RECT 35.800 48.000 36.200 49.900 ;
        RECT 34.200 47.900 36.200 48.000 ;
        RECT 36.600 47.900 37.000 49.900 ;
        RECT 37.700 48.200 38.100 49.900 ;
        RECT 37.700 47.900 38.600 48.200 ;
        RECT 34.300 47.700 36.100 47.900 ;
        RECT 31.900 47.400 33.800 47.700 ;
        RECT 27.800 47.100 28.200 47.200 ;
        RECT 29.900 47.100 30.300 47.200 ;
        RECT 25.000 46.800 30.500 47.100 ;
        RECT 26.500 46.700 26.900 46.800 ;
        RECT 21.400 45.800 23.400 46.100 ;
        RECT 25.700 46.200 26.100 46.300 ;
        RECT 27.000 46.200 27.400 46.300 ;
        RECT 25.700 45.900 28.200 46.200 ;
        RECT 27.800 45.800 28.200 45.900 ;
        RECT 21.400 45.200 21.700 45.800 ;
        RECT 21.400 45.100 21.800 45.200 ;
        RECT 15.800 44.800 16.500 45.100 ;
        RECT 16.800 44.800 17.300 45.100 ;
        RECT 16.200 44.200 16.500 44.800 ;
        RECT 16.200 43.800 16.600 44.200 ;
        RECT 16.900 41.100 17.300 44.800 ;
        RECT 20.300 44.800 20.800 45.100 ;
        RECT 21.100 44.800 21.800 45.100 ;
        RECT 20.300 41.100 20.700 44.800 ;
        RECT 21.100 44.200 21.400 44.800 ;
        RECT 22.200 44.400 22.600 45.200 ;
        RECT 21.000 43.800 21.400 44.200 ;
        RECT 23.000 41.100 23.400 45.800 ;
        RECT 24.600 45.500 27.400 45.600 ;
        RECT 24.600 45.400 27.500 45.500 ;
        RECT 24.600 45.300 29.500 45.400 ;
        RECT 24.600 41.100 25.000 45.300 ;
        RECT 27.100 45.100 29.500 45.300 ;
        RECT 26.200 44.500 28.900 44.800 ;
        RECT 26.200 44.400 26.600 44.500 ;
        RECT 28.500 44.400 28.900 44.500 ;
        RECT 29.200 44.500 29.500 45.100 ;
        RECT 30.200 45.200 30.500 46.800 ;
        RECT 31.000 46.400 31.400 46.500 ;
        RECT 31.000 46.100 32.900 46.400 ;
        RECT 32.500 46.000 32.900 46.100 ;
        RECT 31.700 45.700 32.100 45.800 ;
        RECT 33.400 45.700 33.800 47.400 ;
        RECT 34.600 47.200 35.000 47.400 ;
        RECT 36.600 47.200 36.900 47.900 ;
        RECT 34.200 46.900 35.000 47.200 ;
        RECT 34.200 46.800 34.600 46.900 ;
        RECT 35.700 46.800 37.000 47.200 ;
        RECT 35.000 45.800 35.400 46.600 ;
        RECT 31.700 45.400 33.800 45.700 ;
        RECT 30.200 44.900 31.400 45.200 ;
        RECT 29.900 44.500 30.300 44.600 ;
        RECT 29.200 44.200 30.300 44.500 ;
        RECT 31.100 44.400 31.400 44.900 ;
        RECT 31.100 44.000 31.800 44.400 ;
        RECT 27.900 43.700 28.300 43.800 ;
        RECT 29.300 43.700 29.700 43.800 ;
        RECT 26.200 43.100 26.600 43.500 ;
        RECT 27.900 43.400 29.700 43.700 ;
        RECT 29.000 43.100 29.300 43.400 ;
        RECT 31.000 43.100 31.400 43.500 ;
        RECT 26.200 42.800 27.200 43.100 ;
        RECT 26.800 41.100 27.200 42.800 ;
        RECT 29.000 41.100 29.400 43.100 ;
        RECT 31.100 41.100 31.700 43.100 ;
        RECT 33.400 41.100 33.800 45.400 ;
        RECT 35.700 45.100 36.000 46.800 ;
        RECT 38.200 46.100 38.600 47.900 ;
        RECT 39.000 46.800 39.400 47.600 ;
        RECT 39.800 47.500 40.200 49.900 ;
        RECT 42.000 49.200 42.400 49.900 ;
        RECT 41.400 48.900 42.400 49.200 ;
        RECT 44.200 48.900 44.600 49.900 ;
        RECT 46.300 49.200 46.900 49.900 ;
        RECT 46.200 48.900 46.900 49.200 ;
        RECT 41.400 48.500 41.800 48.900 ;
        RECT 44.200 48.600 44.500 48.900 ;
        RECT 42.200 48.200 42.600 48.600 ;
        RECT 43.100 48.300 44.500 48.600 ;
        RECT 46.200 48.500 46.600 48.900 ;
        RECT 43.100 48.200 43.500 48.300 ;
        RECT 40.200 47.100 41.000 47.200 ;
        RECT 42.300 47.100 42.600 48.200 ;
        RECT 45.400 48.100 45.800 48.200 ;
        RECT 45.400 47.800 47.400 48.100 ;
        RECT 47.000 47.700 47.500 47.800 ;
        RECT 48.600 47.700 49.000 49.900 ;
        RECT 51.000 48.000 51.400 49.900 ;
        RECT 52.600 48.000 53.000 49.900 ;
        RECT 51.000 47.900 53.000 48.000 ;
        RECT 53.400 47.900 53.800 49.900 ;
        RECT 54.200 48.000 54.600 49.900 ;
        RECT 55.800 48.000 56.200 49.900 ;
        RECT 54.200 47.900 56.200 48.000 ;
        RECT 56.600 47.900 57.000 49.900 ;
        RECT 51.100 47.700 52.900 47.900 ;
        RECT 47.000 47.400 49.000 47.700 ;
        RECT 45.100 47.100 45.500 47.200 ;
        RECT 40.200 46.800 45.700 47.100 ;
        RECT 41.700 46.700 42.100 46.800 ;
        RECT 36.600 45.800 38.600 46.100 ;
        RECT 40.900 46.200 41.300 46.300 ;
        RECT 42.200 46.200 42.600 46.300 ;
        RECT 40.900 45.900 43.400 46.200 ;
        RECT 43.000 45.800 43.400 45.900 ;
        RECT 44.600 46.100 45.000 46.200 ;
        RECT 45.400 46.100 45.700 46.800 ;
        RECT 46.200 46.400 46.600 46.500 ;
        RECT 46.200 46.100 48.100 46.400 ;
        RECT 44.600 45.800 45.700 46.100 ;
        RECT 47.700 46.000 48.100 46.100 ;
        RECT 36.600 45.200 36.900 45.800 ;
        RECT 36.600 45.100 37.000 45.200 ;
        RECT 35.500 44.800 36.000 45.100 ;
        RECT 36.300 44.800 37.000 45.100 ;
        RECT 35.500 41.100 35.900 44.800 ;
        RECT 36.300 44.200 36.600 44.800 ;
        RECT 37.400 44.400 37.800 45.200 ;
        RECT 36.200 43.800 36.600 44.200 ;
        RECT 38.200 41.100 38.600 45.800 ;
        RECT 39.800 45.500 42.600 45.600 ;
        RECT 39.800 45.400 42.700 45.500 ;
        RECT 39.800 45.300 44.700 45.400 ;
        RECT 39.800 41.100 40.200 45.300 ;
        RECT 42.300 45.100 44.700 45.300 ;
        RECT 41.400 44.500 44.100 44.800 ;
        RECT 41.400 44.400 41.800 44.500 ;
        RECT 43.700 44.400 44.100 44.500 ;
        RECT 44.400 44.500 44.700 45.100 ;
        RECT 45.400 45.200 45.700 45.800 ;
        RECT 46.900 45.700 47.300 45.800 ;
        RECT 48.600 45.700 49.000 47.400 ;
        RECT 51.400 47.200 51.800 47.400 ;
        RECT 53.400 47.200 53.700 47.900 ;
        RECT 54.300 47.700 56.100 47.900 ;
        RECT 54.600 47.200 55.000 47.400 ;
        RECT 56.600 47.200 56.900 47.900 ;
        RECT 57.400 47.600 57.800 49.900 ;
        RECT 59.000 48.200 59.400 49.900 ;
        RECT 59.000 47.900 59.500 48.200 ;
        RECT 57.400 47.300 58.700 47.600 ;
        RECT 51.000 46.900 51.800 47.200 ;
        RECT 51.000 46.800 51.400 46.900 ;
        RECT 52.500 46.800 53.800 47.200 ;
        RECT 54.200 46.900 55.000 47.200 ;
        RECT 54.200 46.800 54.600 46.900 ;
        RECT 55.700 46.800 57.000 47.200 ;
        RECT 51.800 45.800 52.200 46.600 ;
        RECT 52.500 46.100 52.800 46.800 ;
        RECT 55.000 46.100 55.400 46.600 ;
        RECT 52.500 45.800 55.400 46.100 ;
        RECT 46.900 45.400 49.000 45.700 ;
        RECT 45.400 44.900 46.600 45.200 ;
        RECT 45.100 44.500 45.500 44.600 ;
        RECT 44.400 44.200 45.500 44.500 ;
        RECT 46.300 44.400 46.600 44.900 ;
        RECT 46.300 44.000 47.000 44.400 ;
        RECT 43.100 43.700 43.500 43.800 ;
        RECT 44.500 43.700 44.900 43.800 ;
        RECT 41.400 43.100 41.800 43.500 ;
        RECT 43.100 43.400 44.900 43.700 ;
        RECT 44.200 43.100 44.500 43.400 ;
        RECT 46.200 43.100 46.600 43.500 ;
        RECT 41.400 42.800 42.400 43.100 ;
        RECT 42.000 41.100 42.400 42.800 ;
        RECT 44.200 41.100 44.600 43.100 ;
        RECT 46.300 41.100 46.900 43.100 ;
        RECT 48.600 41.100 49.000 45.400 ;
        RECT 52.500 45.100 52.800 45.800 ;
        RECT 53.400 45.100 53.800 45.200 ;
        RECT 55.700 45.100 56.000 46.800 ;
        RECT 57.500 46.200 57.900 46.600 ;
        RECT 57.400 45.800 57.900 46.200 ;
        RECT 58.400 46.500 58.700 47.300 ;
        RECT 59.200 47.200 59.500 47.900 ;
        RECT 60.600 47.500 61.000 49.900 ;
        RECT 62.800 49.200 63.200 49.900 ;
        RECT 62.200 48.900 63.200 49.200 ;
        RECT 65.000 48.900 65.400 49.900 ;
        RECT 67.100 49.200 67.700 49.900 ;
        RECT 67.000 48.900 67.700 49.200 ;
        RECT 62.200 48.500 62.600 48.900 ;
        RECT 65.000 48.600 65.300 48.900 ;
        RECT 63.000 48.200 63.400 48.600 ;
        RECT 63.900 48.300 65.300 48.600 ;
        RECT 67.000 48.500 67.400 48.900 ;
        RECT 63.900 48.200 64.300 48.300 ;
        RECT 59.000 46.800 59.500 47.200 ;
        RECT 61.000 47.100 61.800 47.200 ;
        RECT 63.100 47.100 63.400 48.200 ;
        RECT 67.900 47.700 68.300 47.800 ;
        RECT 69.400 47.700 69.800 49.900 ;
        RECT 67.900 47.400 69.800 47.700 ;
        RECT 70.200 47.500 70.600 49.900 ;
        RECT 72.400 49.200 72.800 49.900 ;
        RECT 71.800 48.900 72.800 49.200 ;
        RECT 74.600 48.900 75.000 49.900 ;
        RECT 76.700 49.200 77.300 49.900 ;
        RECT 76.600 48.900 77.300 49.200 ;
        RECT 71.800 48.500 72.200 48.900 ;
        RECT 74.600 48.600 74.900 48.900 ;
        RECT 72.600 48.200 73.000 48.600 ;
        RECT 73.500 48.300 74.900 48.600 ;
        RECT 76.600 48.500 77.000 48.900 ;
        RECT 73.500 48.200 73.900 48.300 ;
        RECT 65.900 47.100 66.300 47.200 ;
        RECT 61.000 46.800 66.500 47.100 ;
        RECT 58.400 46.100 58.900 46.500 ;
        RECT 56.600 45.100 57.000 45.200 ;
        RECT 58.400 45.100 58.700 46.100 ;
        RECT 59.200 45.100 59.500 46.800 ;
        RECT 62.500 46.700 62.900 46.800 ;
        RECT 61.700 46.200 62.100 46.300 ;
        RECT 61.700 46.100 64.200 46.200 ;
        RECT 65.400 46.100 65.800 46.200 ;
        RECT 61.700 45.900 65.800 46.100 ;
        RECT 63.800 45.800 65.800 45.900 ;
        RECT 52.300 44.800 52.800 45.100 ;
        RECT 53.100 44.800 53.800 45.100 ;
        RECT 55.500 44.800 56.000 45.100 ;
        RECT 56.300 44.800 57.000 45.100 ;
        RECT 57.400 44.800 58.700 45.100 ;
        RECT 52.300 41.100 52.700 44.800 ;
        RECT 53.100 44.200 53.400 44.800 ;
        RECT 53.000 43.800 53.400 44.200 ;
        RECT 55.500 41.100 55.900 44.800 ;
        RECT 56.300 44.200 56.600 44.800 ;
        RECT 56.200 43.800 56.600 44.200 ;
        RECT 57.400 41.100 57.800 44.800 ;
        RECT 59.000 44.600 59.500 45.100 ;
        RECT 60.600 45.500 63.400 45.600 ;
        RECT 60.600 45.400 63.500 45.500 ;
        RECT 60.600 45.300 65.500 45.400 ;
        RECT 59.000 41.100 59.400 44.600 ;
        RECT 60.600 41.100 61.000 45.300 ;
        RECT 63.100 45.100 65.500 45.300 ;
        RECT 62.200 44.500 64.900 44.800 ;
        RECT 62.200 44.400 62.600 44.500 ;
        RECT 64.500 44.400 64.900 44.500 ;
        RECT 65.200 44.500 65.500 45.100 ;
        RECT 66.200 45.200 66.500 46.800 ;
        RECT 67.000 46.400 67.400 46.500 ;
        RECT 67.000 46.100 68.900 46.400 ;
        RECT 68.500 46.000 68.900 46.100 ;
        RECT 67.700 45.700 68.100 45.800 ;
        RECT 69.400 45.700 69.800 47.400 ;
        RECT 70.600 47.100 71.400 47.200 ;
        RECT 72.700 47.100 73.000 48.200 ;
        RECT 79.000 48.100 79.400 49.900 ;
        RECT 79.800 48.100 80.200 48.600 ;
        RECT 79.000 47.800 80.200 48.100 ;
        RECT 77.500 47.700 77.900 47.800 ;
        RECT 79.000 47.700 79.400 47.800 ;
        RECT 77.500 47.400 79.400 47.700 ;
        RECT 75.500 47.100 75.900 47.200 ;
        RECT 70.600 46.800 76.100 47.100 ;
        RECT 72.100 46.700 72.500 46.800 ;
        RECT 71.300 46.200 71.700 46.300 ;
        RECT 71.300 46.100 73.800 46.200 ;
        RECT 75.000 46.100 75.400 46.200 ;
        RECT 71.300 45.900 75.400 46.100 ;
        RECT 73.400 45.800 75.400 45.900 ;
        RECT 67.700 45.400 69.800 45.700 ;
        RECT 66.200 44.900 67.400 45.200 ;
        RECT 65.900 44.500 66.300 44.600 ;
        RECT 65.200 44.200 66.300 44.500 ;
        RECT 67.100 44.400 67.400 44.900 ;
        RECT 67.100 44.000 67.800 44.400 ;
        RECT 63.900 43.700 64.300 43.800 ;
        RECT 65.300 43.700 65.700 43.800 ;
        RECT 62.200 43.100 62.600 43.500 ;
        RECT 63.900 43.400 65.700 43.700 ;
        RECT 65.000 43.100 65.300 43.400 ;
        RECT 67.000 43.100 67.400 43.500 ;
        RECT 62.200 42.800 63.200 43.100 ;
        RECT 62.800 41.100 63.200 42.800 ;
        RECT 65.000 41.100 65.400 43.100 ;
        RECT 67.100 41.100 67.700 43.100 ;
        RECT 69.400 41.100 69.800 45.400 ;
        RECT 70.200 45.500 73.000 45.600 ;
        RECT 70.200 45.400 73.100 45.500 ;
        RECT 70.200 45.300 75.100 45.400 ;
        RECT 70.200 41.100 70.600 45.300 ;
        RECT 72.700 45.100 75.100 45.300 ;
        RECT 71.800 44.500 74.500 44.800 ;
        RECT 71.800 44.400 72.200 44.500 ;
        RECT 74.100 44.400 74.500 44.500 ;
        RECT 74.800 44.500 75.100 45.100 ;
        RECT 75.800 45.200 76.100 46.800 ;
        RECT 76.600 46.400 77.000 46.500 ;
        RECT 76.600 46.100 78.500 46.400 ;
        RECT 78.100 46.000 78.500 46.100 ;
        RECT 77.300 45.700 77.700 45.800 ;
        RECT 79.000 45.700 79.400 47.400 ;
        RECT 77.300 45.400 79.400 45.700 ;
        RECT 75.800 44.900 77.000 45.200 ;
        RECT 75.500 44.500 75.900 44.600 ;
        RECT 74.800 44.200 75.900 44.500 ;
        RECT 76.700 44.400 77.000 44.900 ;
        RECT 76.700 44.000 77.400 44.400 ;
        RECT 73.500 43.700 73.900 43.800 ;
        RECT 74.900 43.700 75.300 43.800 ;
        RECT 71.800 43.100 72.200 43.500 ;
        RECT 73.500 43.400 75.300 43.700 ;
        RECT 74.600 43.100 74.900 43.400 ;
        RECT 76.600 43.100 77.000 43.500 ;
        RECT 71.800 42.800 72.800 43.100 ;
        RECT 72.400 41.100 72.800 42.800 ;
        RECT 74.600 41.100 75.000 43.100 ;
        RECT 76.700 41.100 77.300 43.100 ;
        RECT 79.000 41.100 79.400 45.400 ;
        RECT 80.600 41.100 81.000 49.900 ;
        RECT 83.300 48.000 83.700 49.500 ;
        RECT 85.400 48.500 85.800 49.500 ;
        RECT 82.900 47.700 83.700 48.000 ;
        RECT 82.900 47.500 83.300 47.700 ;
        RECT 82.900 47.200 83.200 47.500 ;
        RECT 85.500 47.400 85.800 48.500 ;
        RECT 82.200 46.800 83.200 47.200 ;
        RECT 83.700 47.100 85.800 47.400 ;
        RECT 87.000 48.800 87.400 49.900 ;
        RECT 87.000 47.200 87.300 48.800 ;
        RECT 87.800 47.800 88.200 48.600 ;
        RECT 90.200 47.900 90.600 49.900 ;
        RECT 90.900 48.200 91.300 48.600 ;
        RECT 83.700 46.900 84.200 47.100 ;
        RECT 82.200 45.400 82.600 46.200 ;
        RECT 82.900 44.900 83.200 46.800 ;
        RECT 83.500 46.500 84.200 46.900 ;
        RECT 87.000 46.800 87.400 47.200 ;
        RECT 83.900 45.500 84.200 46.500 ;
        RECT 84.600 45.800 85.000 46.600 ;
        RECT 85.400 45.800 85.800 46.600 ;
        RECT 83.900 45.200 85.800 45.500 ;
        RECT 86.200 45.400 86.600 46.200 ;
        RECT 82.900 44.600 83.700 44.900 ;
        RECT 83.300 41.100 83.700 44.600 ;
        RECT 85.500 43.500 85.800 45.200 ;
        RECT 87.000 45.100 87.300 46.800 ;
        RECT 89.400 46.400 89.800 47.200 ;
        RECT 88.600 46.100 89.000 46.200 ;
        RECT 90.200 46.100 90.500 47.900 ;
        RECT 91.000 47.800 91.400 48.200 ;
        RECT 91.800 48.000 92.200 49.900 ;
        RECT 93.400 48.000 93.800 49.900 ;
        RECT 91.800 47.900 93.800 48.000 ;
        RECT 94.200 47.900 94.600 49.900 ;
        RECT 95.000 47.900 95.400 49.900 ;
        RECT 95.800 48.000 96.200 49.900 ;
        RECT 97.400 48.000 97.800 49.900 ;
        RECT 95.800 47.900 97.800 48.000 ;
        RECT 91.900 47.700 93.700 47.900 ;
        RECT 92.200 47.200 92.600 47.400 ;
        RECT 94.200 47.200 94.500 47.900 ;
        RECT 95.100 47.200 95.400 47.900 ;
        RECT 95.900 47.700 97.700 47.900 ;
        RECT 98.200 47.600 98.600 49.900 ;
        RECT 99.800 48.200 100.200 49.900 ;
        RECT 99.800 47.900 100.300 48.200 ;
        RECT 97.000 47.200 97.400 47.400 ;
        RECT 98.200 47.300 99.500 47.600 ;
        RECT 91.800 46.900 92.600 47.200 ;
        RECT 91.800 46.800 92.200 46.900 ;
        RECT 93.300 46.800 94.600 47.200 ;
        RECT 95.000 46.800 96.300 47.200 ;
        RECT 97.000 46.900 97.800 47.200 ;
        RECT 97.400 46.800 97.800 46.900 ;
        RECT 91.000 46.100 91.400 46.200 ;
        RECT 88.600 45.800 89.400 46.100 ;
        RECT 90.200 45.800 91.400 46.100 ;
        RECT 92.600 45.800 93.000 46.600 ;
        RECT 89.000 45.600 89.400 45.800 ;
        RECT 91.000 45.100 91.300 45.800 ;
        RECT 93.300 45.100 93.600 46.800 ;
        RECT 94.200 45.100 94.600 45.200 ;
        RECT 85.400 41.500 85.800 43.500 ;
        RECT 86.500 44.700 87.400 45.100 ;
        RECT 88.600 44.800 90.600 45.100 ;
        RECT 86.500 41.100 86.900 44.700 ;
        RECT 88.600 41.100 89.000 44.800 ;
        RECT 90.200 41.100 90.600 44.800 ;
        RECT 91.000 41.100 91.400 45.100 ;
        RECT 93.100 44.800 93.600 45.100 ;
        RECT 93.900 44.800 94.600 45.100 ;
        RECT 95.000 45.100 95.400 45.200 ;
        RECT 96.000 45.100 96.300 46.800 ;
        RECT 96.600 45.800 97.000 46.600 ;
        RECT 98.300 46.200 98.700 46.600 ;
        RECT 98.200 45.800 98.700 46.200 ;
        RECT 99.200 46.500 99.500 47.300 ;
        RECT 100.000 47.200 100.300 47.900 ;
        RECT 104.600 47.900 105.000 49.900 ;
        RECT 105.300 48.200 105.700 48.600 ;
        RECT 99.800 47.100 100.300 47.200 ;
        RECT 100.600 47.100 101.000 47.200 ;
        RECT 99.800 46.800 101.000 47.100 ;
        RECT 99.200 46.100 99.700 46.500 ;
        RECT 99.200 45.100 99.500 46.100 ;
        RECT 100.000 45.100 100.300 46.800 ;
        RECT 103.800 46.400 104.200 47.200 ;
        RECT 103.000 46.100 103.400 46.200 ;
        RECT 104.600 46.100 104.900 47.900 ;
        RECT 105.400 47.800 105.800 48.200 ;
        RECT 107.800 47.900 108.200 49.900 ;
        RECT 108.500 48.200 108.900 48.600 ;
        RECT 109.500 48.200 109.900 48.600 ;
        RECT 107.000 46.400 107.400 47.200 ;
        RECT 105.400 46.100 105.800 46.200 ;
        RECT 103.000 45.800 103.800 46.100 ;
        RECT 104.600 45.800 105.800 46.100 ;
        RECT 106.200 46.100 106.600 46.200 ;
        RECT 107.800 46.100 108.100 47.900 ;
        RECT 108.600 47.800 109.000 48.200 ;
        RECT 109.400 47.800 109.800 48.200 ;
        RECT 110.200 47.900 110.600 49.900 ;
        RECT 112.600 47.900 113.000 49.900 ;
        RECT 113.400 48.000 113.800 49.900 ;
        RECT 115.000 48.000 115.400 49.900 ;
        RECT 113.400 47.900 115.400 48.000 ;
        RECT 116.600 48.800 117.000 49.900 ;
        RECT 108.600 46.100 109.000 46.200 ;
        RECT 106.200 45.800 107.000 46.100 ;
        RECT 107.800 45.800 109.000 46.100 ;
        RECT 109.400 46.100 109.800 46.200 ;
        RECT 110.300 46.100 110.600 47.900 ;
        RECT 112.700 47.200 113.000 47.900 ;
        RECT 113.500 47.700 115.300 47.900 ;
        RECT 114.600 47.200 115.000 47.400 ;
        RECT 116.600 47.200 116.900 48.800 ;
        RECT 117.400 48.100 117.800 48.600 ;
        RECT 118.200 48.100 118.600 49.900 ;
        RECT 120.300 49.200 120.900 49.900 ;
        RECT 120.300 48.900 121.000 49.200 ;
        RECT 122.600 48.900 123.000 49.900 ;
        RECT 124.800 49.200 125.200 49.900 ;
        RECT 124.800 48.900 125.800 49.200 ;
        RECT 120.600 48.500 121.000 48.900 ;
        RECT 122.700 48.600 123.000 48.900 ;
        RECT 122.700 48.300 124.100 48.600 ;
        RECT 123.700 48.200 124.100 48.300 ;
        RECT 117.400 47.800 118.600 48.100 ;
        RECT 124.600 47.800 125.000 48.600 ;
        RECT 125.400 48.500 125.800 48.900 ;
        RECT 118.200 47.700 118.600 47.800 ;
        RECT 119.700 47.700 120.100 47.800 ;
        RECT 118.200 47.400 120.100 47.700 ;
        RECT 111.000 46.400 111.400 47.200 ;
        RECT 111.800 47.100 112.200 47.200 ;
        RECT 112.600 47.100 113.900 47.200 ;
        RECT 111.800 46.800 113.900 47.100 ;
        RECT 114.600 46.900 115.400 47.200 ;
        RECT 115.000 46.800 115.400 46.900 ;
        RECT 116.600 46.800 117.000 47.200 ;
        RECT 111.800 46.100 112.200 46.200 ;
        RECT 109.400 45.800 110.600 46.100 ;
        RECT 111.400 45.800 112.200 46.100 ;
        RECT 103.400 45.600 103.800 45.800 ;
        RECT 105.400 45.100 105.700 45.800 ;
        RECT 106.600 45.600 107.000 45.800 ;
        RECT 108.600 45.100 108.900 45.800 ;
        RECT 109.500 45.100 109.800 45.800 ;
        RECT 111.400 45.600 111.800 45.800 ;
        RECT 112.600 45.100 113.000 45.200 ;
        RECT 113.600 45.100 113.900 46.800 ;
        RECT 114.200 45.800 114.600 46.600 ;
        RECT 115.800 45.400 116.200 46.200 ;
        RECT 116.600 45.100 116.900 46.800 ;
        RECT 118.200 45.700 118.600 47.400 ;
        RECT 121.700 47.100 122.100 47.200 ;
        RECT 124.600 47.100 124.900 47.800 ;
        RECT 127.000 47.500 127.400 49.900 ;
        RECT 127.800 47.900 128.200 49.900 ;
        RECT 128.600 48.000 129.000 49.900 ;
        RECT 130.200 48.000 130.600 49.900 ;
        RECT 131.800 48.200 132.200 49.900 ;
        RECT 128.600 47.900 130.600 48.000 ;
        RECT 131.700 47.900 132.200 48.200 ;
        RECT 127.900 47.200 128.200 47.900 ;
        RECT 128.700 47.700 130.500 47.900 ;
        RECT 129.800 47.200 130.200 47.400 ;
        RECT 131.700 47.200 132.000 47.900 ;
        RECT 133.400 47.600 133.800 49.900 ;
        RECT 132.500 47.300 133.800 47.600 ;
        RECT 134.200 47.700 134.600 49.900 ;
        RECT 136.300 49.200 136.900 49.900 ;
        RECT 136.300 48.900 137.000 49.200 ;
        RECT 138.600 48.900 139.000 49.900 ;
        RECT 140.800 49.200 141.200 49.900 ;
        RECT 140.800 48.900 141.800 49.200 ;
        RECT 136.600 48.500 137.000 48.900 ;
        RECT 138.700 48.600 139.000 48.900 ;
        RECT 138.700 48.300 140.100 48.600 ;
        RECT 139.700 48.200 140.100 48.300 ;
        RECT 140.600 48.200 141.000 48.600 ;
        RECT 141.400 48.500 141.800 48.900 ;
        RECT 135.700 47.700 136.100 47.800 ;
        RECT 134.200 47.400 136.100 47.700 ;
        RECT 126.200 47.100 127.000 47.200 ;
        RECT 121.500 46.800 127.000 47.100 ;
        RECT 127.800 46.800 129.100 47.200 ;
        RECT 129.800 47.100 130.600 47.200 ;
        RECT 131.700 47.100 132.200 47.200 ;
        RECT 129.800 46.900 132.200 47.100 ;
        RECT 130.200 46.800 132.200 46.900 ;
        RECT 120.600 46.400 121.000 46.500 ;
        RECT 119.100 46.100 121.000 46.400 ;
        RECT 119.100 46.000 119.500 46.100 ;
        RECT 119.900 45.700 120.300 45.800 ;
        RECT 118.200 45.400 120.300 45.700 ;
        RECT 95.000 44.800 95.700 45.100 ;
        RECT 96.000 44.800 96.500 45.100 ;
        RECT 93.100 41.100 93.500 44.800 ;
        RECT 93.900 44.200 94.200 44.800 ;
        RECT 93.800 43.800 94.200 44.200 ;
        RECT 95.400 44.200 95.700 44.800 ;
        RECT 95.400 43.800 95.800 44.200 ;
        RECT 96.100 41.100 96.500 44.800 ;
        RECT 98.200 44.800 99.500 45.100 ;
        RECT 98.200 41.100 98.600 44.800 ;
        RECT 99.800 44.600 100.300 45.100 ;
        RECT 103.000 44.800 105.000 45.100 ;
        RECT 99.800 41.100 100.200 44.600 ;
        RECT 103.000 41.100 103.400 44.800 ;
        RECT 104.600 41.100 105.000 44.800 ;
        RECT 105.400 41.100 105.800 45.100 ;
        RECT 106.200 44.800 108.200 45.100 ;
        RECT 106.200 41.100 106.600 44.800 ;
        RECT 107.800 41.100 108.200 44.800 ;
        RECT 108.600 41.100 109.000 45.100 ;
        RECT 109.400 41.100 109.800 45.100 ;
        RECT 110.200 44.800 112.200 45.100 ;
        RECT 112.600 44.800 113.300 45.100 ;
        RECT 113.600 44.800 114.100 45.100 ;
        RECT 110.200 41.100 110.600 44.800 ;
        RECT 111.800 41.100 112.200 44.800 ;
        RECT 113.000 44.200 113.300 44.800 ;
        RECT 113.000 43.800 113.400 44.200 ;
        RECT 113.700 41.100 114.100 44.800 ;
        RECT 116.100 44.700 117.000 45.100 ;
        RECT 116.100 41.100 116.500 44.700 ;
        RECT 118.200 41.100 118.600 45.400 ;
        RECT 121.500 45.200 121.800 46.800 ;
        RECT 125.100 46.700 125.500 46.800 ;
        RECT 125.900 46.200 126.300 46.300 ;
        RECT 122.200 46.100 122.600 46.200 ;
        RECT 123.800 46.100 126.300 46.200 ;
        RECT 122.200 45.900 126.300 46.100 ;
        RECT 127.800 46.200 128.100 46.800 ;
        RECT 122.200 45.800 124.200 45.900 ;
        RECT 127.800 45.800 128.200 46.200 ;
        RECT 124.600 45.500 127.400 45.600 ;
        RECT 124.500 45.400 127.400 45.500 ;
        RECT 120.600 44.900 121.800 45.200 ;
        RECT 122.500 45.300 127.400 45.400 ;
        RECT 122.500 45.100 124.900 45.300 ;
        RECT 120.600 44.400 120.900 44.900 ;
        RECT 120.200 44.000 120.900 44.400 ;
        RECT 121.700 44.500 122.100 44.600 ;
        RECT 122.500 44.500 122.800 45.100 ;
        RECT 121.700 44.200 122.800 44.500 ;
        RECT 123.100 44.500 125.800 44.800 ;
        RECT 123.100 44.400 123.500 44.500 ;
        RECT 125.400 44.400 125.800 44.500 ;
        RECT 122.300 43.700 122.700 43.800 ;
        RECT 123.700 43.700 124.100 43.800 ;
        RECT 120.600 43.100 121.000 43.500 ;
        RECT 122.300 43.400 124.100 43.700 ;
        RECT 122.700 43.100 123.000 43.400 ;
        RECT 125.400 43.100 125.800 43.500 ;
        RECT 120.300 41.100 120.900 43.100 ;
        RECT 122.600 41.100 123.000 43.100 ;
        RECT 124.800 42.800 125.800 43.100 ;
        RECT 124.800 41.100 125.200 42.800 ;
        RECT 127.000 41.100 127.400 45.300 ;
        RECT 127.800 45.100 128.200 45.200 ;
        RECT 128.800 45.100 129.100 46.800 ;
        RECT 129.400 45.800 129.800 46.600 ;
        RECT 131.700 45.100 132.000 46.800 ;
        RECT 132.500 46.500 132.800 47.300 ;
        RECT 132.300 46.100 132.800 46.500 ;
        RECT 132.500 45.100 132.800 46.100 ;
        RECT 133.300 46.200 133.700 46.600 ;
        RECT 133.300 45.800 133.800 46.200 ;
        RECT 134.200 45.700 134.600 47.400 ;
        RECT 137.700 47.100 138.100 47.200 ;
        RECT 139.800 47.100 140.200 47.200 ;
        RECT 140.600 47.100 140.900 48.200 ;
        RECT 143.000 47.500 143.400 49.900 ;
        RECT 144.600 48.900 145.000 49.900 ;
        RECT 143.800 47.800 144.200 48.600 ;
        RECT 144.700 48.100 145.000 48.900 ;
        RECT 146.300 48.200 146.700 48.600 ;
        RECT 146.200 48.100 146.600 48.200 ;
        RECT 144.600 47.800 146.600 48.100 ;
        RECT 147.000 47.900 147.400 49.900 ;
        RECT 144.700 47.200 145.000 47.800 ;
        RECT 142.200 47.100 143.000 47.200 ;
        RECT 137.500 46.800 143.000 47.100 ;
        RECT 144.600 46.800 145.000 47.200 ;
        RECT 136.600 46.400 137.000 46.500 ;
        RECT 135.100 46.100 137.000 46.400 ;
        RECT 135.100 46.000 135.500 46.100 ;
        RECT 135.900 45.700 136.300 45.800 ;
        RECT 134.200 45.400 136.300 45.700 ;
        RECT 127.800 44.800 128.500 45.100 ;
        RECT 128.800 44.800 129.300 45.100 ;
        RECT 128.200 44.200 128.500 44.800 ;
        RECT 128.200 43.800 128.600 44.200 ;
        RECT 128.900 41.100 129.300 44.800 ;
        RECT 131.700 44.600 132.200 45.100 ;
        RECT 132.500 44.800 133.800 45.100 ;
        RECT 131.800 41.100 132.200 44.600 ;
        RECT 133.400 41.100 133.800 44.800 ;
        RECT 134.200 41.100 134.600 45.400 ;
        RECT 137.500 45.200 137.800 46.800 ;
        RECT 141.100 46.700 141.500 46.800 ;
        RECT 140.600 46.200 141.000 46.300 ;
        RECT 141.900 46.200 142.300 46.300 ;
        RECT 139.800 45.900 142.300 46.200 ;
        RECT 139.800 45.800 140.200 45.900 ;
        RECT 140.600 45.500 143.400 45.600 ;
        RECT 140.500 45.400 143.400 45.500 ;
        RECT 136.600 44.900 137.800 45.200 ;
        RECT 138.500 45.300 143.400 45.400 ;
        RECT 138.500 45.100 140.900 45.300 ;
        RECT 136.600 44.400 136.900 44.900 ;
        RECT 136.200 44.000 136.900 44.400 ;
        RECT 137.700 44.500 138.100 44.600 ;
        RECT 138.500 44.500 138.800 45.100 ;
        RECT 137.700 44.200 138.800 44.500 ;
        RECT 139.100 44.500 141.800 44.800 ;
        RECT 139.100 44.400 139.500 44.500 ;
        RECT 141.400 44.400 141.800 44.500 ;
        RECT 138.300 43.700 138.700 43.800 ;
        RECT 139.700 43.700 140.100 43.800 ;
        RECT 136.600 43.100 137.000 43.500 ;
        RECT 138.300 43.400 140.100 43.700 ;
        RECT 138.700 43.100 139.000 43.400 ;
        RECT 141.400 43.100 141.800 43.500 ;
        RECT 136.300 41.100 136.900 43.100 ;
        RECT 138.600 41.100 139.000 43.100 ;
        RECT 140.800 42.800 141.800 43.100 ;
        RECT 140.800 41.100 141.200 42.800 ;
        RECT 143.000 41.100 143.400 45.300 ;
        RECT 144.700 45.100 145.000 46.800 ;
        RECT 146.200 46.800 146.600 47.200 ;
        RECT 146.200 46.200 146.500 46.800 ;
        RECT 145.400 45.400 145.800 46.200 ;
        RECT 146.200 46.100 146.600 46.200 ;
        RECT 147.100 46.100 147.400 47.900 ;
        RECT 149.400 47.800 149.800 49.900 ;
        RECT 150.200 48.000 150.600 49.900 ;
        RECT 151.800 48.000 152.200 49.900 ;
        RECT 150.200 47.900 152.200 48.000 ;
        RECT 149.500 47.200 149.800 47.800 ;
        RECT 150.300 47.700 152.100 47.900 ;
        RECT 151.400 47.200 151.800 47.400 ;
        RECT 147.800 46.400 148.200 47.200 ;
        RECT 149.400 46.800 150.700 47.200 ;
        RECT 151.400 46.900 152.200 47.200 ;
        RECT 151.800 46.800 152.200 46.900 ;
        RECT 148.600 46.100 149.000 46.200 ;
        RECT 146.200 45.800 147.400 46.100 ;
        RECT 148.200 45.800 149.000 46.100 ;
        RECT 146.300 45.100 146.600 45.800 ;
        RECT 148.200 45.600 148.600 45.800 ;
        RECT 149.400 45.100 149.800 45.200 ;
        RECT 150.400 45.100 150.700 46.800 ;
        RECT 151.000 45.800 151.400 46.600 ;
        RECT 144.600 44.700 145.500 45.100 ;
        RECT 145.100 41.100 145.500 44.700 ;
        RECT 146.200 41.100 146.600 45.100 ;
        RECT 147.000 44.800 149.000 45.100 ;
        RECT 149.400 44.800 150.100 45.100 ;
        RECT 150.400 44.800 150.900 45.100 ;
        RECT 147.000 41.100 147.400 44.800 ;
        RECT 148.600 41.100 149.000 44.800 ;
        RECT 149.800 44.200 150.100 44.800 ;
        RECT 149.800 43.800 150.200 44.200 ;
        RECT 150.500 41.100 150.900 44.800 ;
        RECT 155.000 41.100 155.400 49.900 ;
        RECT 156.600 48.500 157.000 49.500 ;
        RECT 156.600 47.400 156.900 48.500 ;
        RECT 158.700 48.000 159.100 49.500 ;
        RECT 158.700 47.700 159.500 48.000 ;
        RECT 159.100 47.500 159.500 47.700 ;
        RECT 156.600 47.100 158.700 47.400 ;
        RECT 158.200 46.900 158.700 47.100 ;
        RECT 159.200 47.200 159.500 47.500 ;
        RECT 163.000 47.900 163.400 49.900 ;
        RECT 163.700 48.200 164.100 48.600 ;
        RECT 163.800 48.100 164.200 48.200 ;
        RECT 164.600 48.100 165.000 49.900 ;
        RECT 155.800 46.100 156.200 46.200 ;
        RECT 156.600 46.100 157.000 46.600 ;
        RECT 155.800 45.800 157.000 46.100 ;
        RECT 157.400 45.800 157.800 46.600 ;
        RECT 158.200 46.500 158.900 46.900 ;
        RECT 159.200 46.800 160.200 47.200 ;
        RECT 158.200 45.500 158.500 46.500 ;
        RECT 156.600 45.200 158.500 45.500 ;
        RECT 156.600 43.500 156.900 45.200 ;
        RECT 159.200 44.900 159.500 46.800 ;
        RECT 162.200 46.400 162.600 47.200 ;
        RECT 159.800 45.400 160.200 46.200 ;
        RECT 161.400 46.100 161.800 46.200 ;
        RECT 163.000 46.100 163.300 47.900 ;
        RECT 163.800 47.800 165.000 48.100 ;
        RECT 165.400 48.000 165.800 49.900 ;
        RECT 167.000 48.000 167.400 49.900 ;
        RECT 169.100 48.200 169.500 49.900 ;
        RECT 165.400 47.900 167.400 48.000 ;
        RECT 168.600 47.900 169.500 48.200 ;
        RECT 170.500 48.200 170.900 49.900 ;
        RECT 170.500 47.900 171.400 48.200 ;
        RECT 164.700 47.200 165.000 47.800 ;
        RECT 165.500 47.700 167.300 47.900 ;
        RECT 166.600 47.200 167.000 47.400 ;
        RECT 164.600 46.800 165.900 47.200 ;
        RECT 166.600 46.900 167.400 47.200 ;
        RECT 167.000 46.800 167.400 46.900 ;
        RECT 163.800 46.100 164.200 46.200 ;
        RECT 161.400 45.800 162.200 46.100 ;
        RECT 163.000 45.800 164.200 46.100 ;
        RECT 161.800 45.600 162.200 45.800 ;
        RECT 163.800 45.100 164.100 45.800 ;
        RECT 164.600 45.100 165.000 45.200 ;
        RECT 165.600 45.100 165.900 46.800 ;
        RECT 166.200 46.100 166.600 46.600 ;
        RECT 167.000 46.100 167.400 46.200 ;
        RECT 166.200 45.800 167.400 46.100 ;
        RECT 158.700 44.600 159.500 44.900 ;
        RECT 161.400 44.800 163.400 45.100 ;
        RECT 156.600 41.500 157.000 43.500 ;
        RECT 158.700 42.200 159.100 44.600 ;
        RECT 158.700 41.800 159.400 42.200 ;
        RECT 158.700 41.100 159.100 41.800 ;
        RECT 161.400 41.100 161.800 44.800 ;
        RECT 163.000 41.100 163.400 44.800 ;
        RECT 163.800 41.100 164.200 45.100 ;
        RECT 164.600 44.800 165.300 45.100 ;
        RECT 165.600 44.800 166.100 45.100 ;
        RECT 165.000 44.200 165.300 44.800 ;
        RECT 165.000 43.800 165.400 44.200 ;
        RECT 165.700 41.100 166.100 44.800 ;
        RECT 168.600 41.100 169.000 47.900 ;
        RECT 169.400 45.100 169.800 45.200 ;
        RECT 170.200 45.100 170.600 45.200 ;
        RECT 169.400 44.800 170.600 45.100 ;
        RECT 169.400 44.400 169.800 44.800 ;
        RECT 170.200 44.400 170.600 44.800 ;
        RECT 171.000 41.100 171.400 47.900 ;
        RECT 173.400 41.100 173.800 49.900 ;
        RECT 175.000 47.500 175.400 49.900 ;
        RECT 177.200 49.200 177.600 49.900 ;
        RECT 176.600 48.900 177.600 49.200 ;
        RECT 179.400 48.900 179.800 49.900 ;
        RECT 181.500 49.200 182.100 49.900 ;
        RECT 181.400 48.900 182.100 49.200 ;
        RECT 176.600 48.500 177.000 48.900 ;
        RECT 179.400 48.600 179.700 48.900 ;
        RECT 177.400 48.200 177.800 48.600 ;
        RECT 178.300 48.300 179.700 48.600 ;
        RECT 181.400 48.500 181.800 48.900 ;
        RECT 178.300 48.200 178.700 48.300 ;
        RECT 175.400 47.100 176.200 47.200 ;
        RECT 177.500 47.100 177.800 48.200 ;
        RECT 183.800 48.100 184.200 49.900 ;
        RECT 184.600 48.100 185.000 48.600 ;
        RECT 183.800 47.800 185.000 48.100 ;
        RECT 182.300 47.700 182.700 47.800 ;
        RECT 183.800 47.700 184.200 47.800 ;
        RECT 182.300 47.400 184.200 47.700 ;
        RECT 180.300 47.100 180.700 47.200 ;
        RECT 175.400 46.800 180.900 47.100 ;
        RECT 176.900 46.700 177.300 46.800 ;
        RECT 176.100 46.200 176.500 46.300 ;
        RECT 180.600 46.200 180.900 46.800 ;
        RECT 181.400 46.400 181.800 46.500 ;
        RECT 176.100 45.900 178.600 46.200 ;
        RECT 178.200 45.800 178.600 45.900 ;
        RECT 180.600 45.800 181.000 46.200 ;
        RECT 181.400 46.100 183.300 46.400 ;
        RECT 182.900 46.000 183.300 46.100 ;
        RECT 175.000 45.500 177.800 45.600 ;
        RECT 175.000 45.400 177.900 45.500 ;
        RECT 175.000 45.300 179.900 45.400 ;
        RECT 175.000 41.100 175.400 45.300 ;
        RECT 177.500 45.100 179.900 45.300 ;
        RECT 176.600 44.500 179.300 44.800 ;
        RECT 176.600 44.400 177.000 44.500 ;
        RECT 178.900 44.400 179.300 44.500 ;
        RECT 179.600 44.500 179.900 45.100 ;
        RECT 180.600 45.200 180.900 45.800 ;
        RECT 182.100 45.700 182.500 45.800 ;
        RECT 183.800 45.700 184.200 47.400 ;
        RECT 182.100 45.400 184.200 45.700 ;
        RECT 180.600 44.900 181.800 45.200 ;
        RECT 180.300 44.500 180.700 44.600 ;
        RECT 179.600 44.200 180.700 44.500 ;
        RECT 181.500 44.400 181.800 44.900 ;
        RECT 181.500 44.000 182.200 44.400 ;
        RECT 178.300 43.700 178.700 43.800 ;
        RECT 179.700 43.700 180.100 43.800 ;
        RECT 176.600 43.100 177.000 43.500 ;
        RECT 178.300 43.400 180.100 43.700 ;
        RECT 179.400 43.100 179.700 43.400 ;
        RECT 181.400 43.100 181.800 43.500 ;
        RECT 176.600 42.800 177.600 43.100 ;
        RECT 177.200 41.100 177.600 42.800 ;
        RECT 179.400 41.100 179.800 43.100 ;
        RECT 181.500 41.100 182.100 43.100 ;
        RECT 183.800 41.100 184.200 45.400 ;
        RECT 185.400 41.100 185.800 49.900 ;
        RECT 186.200 48.500 186.600 49.500 ;
        RECT 186.200 47.400 186.500 48.500 ;
        RECT 188.300 48.200 188.700 49.500 ;
        RECT 187.800 48.000 188.700 48.200 ;
        RECT 187.800 47.800 189.100 48.000 ;
        RECT 188.300 47.700 189.100 47.800 ;
        RECT 188.700 47.500 189.100 47.700 ;
        RECT 191.000 47.500 191.400 49.900 ;
        RECT 193.200 49.200 193.600 49.900 ;
        RECT 192.600 48.900 193.600 49.200 ;
        RECT 195.400 48.900 195.800 49.900 ;
        RECT 197.500 49.200 198.100 49.900 ;
        RECT 197.400 48.900 198.100 49.200 ;
        RECT 192.600 48.500 193.000 48.900 ;
        RECT 195.400 48.600 195.700 48.900 ;
        RECT 193.400 48.200 193.800 48.600 ;
        RECT 194.300 48.300 195.700 48.600 ;
        RECT 197.400 48.500 197.800 48.900 ;
        RECT 194.300 48.200 194.700 48.300 ;
        RECT 186.200 47.100 188.300 47.400 ;
        RECT 187.800 46.900 188.300 47.100 ;
        RECT 188.800 47.200 189.100 47.500 ;
        RECT 186.200 45.800 186.600 46.600 ;
        RECT 187.000 45.800 187.400 46.600 ;
        RECT 187.800 46.500 188.500 46.900 ;
        RECT 188.800 46.800 189.800 47.200 ;
        RECT 191.400 47.100 192.200 47.200 ;
        RECT 193.500 47.100 193.800 48.200 ;
        RECT 198.300 47.700 198.700 47.800 ;
        RECT 199.800 47.700 200.200 49.900 ;
        RECT 198.300 47.400 200.200 47.700 ;
        RECT 196.300 47.100 196.700 47.200 ;
        RECT 191.400 46.800 196.900 47.100 ;
        RECT 199.000 46.800 199.400 47.400 ;
        RECT 187.800 45.500 188.100 46.500 ;
        RECT 186.200 45.200 188.100 45.500 ;
        RECT 186.200 43.500 186.500 45.200 ;
        RECT 188.800 44.900 189.100 46.800 ;
        RECT 192.900 46.700 193.300 46.800 ;
        RECT 192.100 46.200 192.500 46.300 ;
        RECT 189.400 46.100 189.800 46.200 ;
        RECT 190.200 46.100 190.600 46.200 ;
        RECT 189.400 45.800 190.600 46.100 ;
        RECT 192.100 46.100 194.600 46.200 ;
        RECT 195.800 46.100 196.200 46.200 ;
        RECT 192.100 45.900 196.200 46.100 ;
        RECT 194.200 45.800 196.200 45.900 ;
        RECT 189.400 45.400 189.800 45.800 ;
        RECT 191.000 45.500 193.800 45.600 ;
        RECT 191.000 45.400 193.900 45.500 ;
        RECT 188.300 44.600 189.100 44.900 ;
        RECT 191.000 45.300 195.900 45.400 ;
        RECT 186.200 41.500 186.600 43.500 ;
        RECT 188.300 41.100 188.700 44.600 ;
        RECT 191.000 41.100 191.400 45.300 ;
        RECT 193.500 45.100 195.900 45.300 ;
        RECT 192.600 44.500 195.300 44.800 ;
        RECT 192.600 44.400 193.000 44.500 ;
        RECT 194.900 44.400 195.300 44.500 ;
        RECT 195.600 44.500 195.900 45.100 ;
        RECT 196.600 45.200 196.900 46.800 ;
        RECT 197.400 46.400 197.800 46.500 ;
        RECT 197.400 46.100 199.300 46.400 ;
        RECT 198.900 46.000 199.300 46.100 ;
        RECT 198.100 45.700 198.500 45.800 ;
        RECT 199.800 45.700 200.200 47.400 ;
        RECT 198.100 45.400 200.200 45.700 ;
        RECT 196.600 44.900 197.800 45.200 ;
        RECT 196.300 44.500 196.700 44.600 ;
        RECT 195.600 44.200 196.700 44.500 ;
        RECT 197.500 44.400 197.800 44.900 ;
        RECT 197.500 44.200 198.200 44.400 ;
        RECT 197.500 44.000 198.600 44.200 ;
        RECT 197.900 43.800 198.600 44.000 ;
        RECT 194.300 43.700 194.700 43.800 ;
        RECT 195.700 43.700 196.100 43.800 ;
        RECT 192.600 43.100 193.000 43.500 ;
        RECT 194.300 43.400 196.100 43.700 ;
        RECT 195.400 43.100 195.700 43.400 ;
        RECT 197.400 43.100 197.800 43.500 ;
        RECT 192.600 42.800 193.600 43.100 ;
        RECT 193.200 41.100 193.600 42.800 ;
        RECT 195.400 41.100 195.800 43.100 ;
        RECT 197.500 41.100 198.100 43.100 ;
        RECT 199.800 41.100 200.200 45.400 ;
        RECT 201.400 41.100 201.800 49.900 ;
        RECT 203.800 48.900 204.200 49.900 ;
        RECT 203.000 47.800 203.400 48.600 ;
        RECT 203.900 47.200 204.200 48.900 ;
        RECT 202.200 47.100 202.600 47.200 ;
        RECT 203.800 47.100 204.200 47.200 ;
        RECT 202.200 46.800 204.200 47.100 ;
        RECT 203.900 45.100 204.200 46.800 ;
        RECT 204.600 45.400 205.000 46.200 ;
        RECT 203.800 44.700 204.700 45.100 ;
        RECT 204.300 41.100 204.700 44.700 ;
        RECT 0.600 35.100 1.000 35.200 ;
        RECT 1.400 35.100 1.800 39.900 ;
        RECT 2.200 35.700 2.600 39.900 ;
        RECT 4.400 38.200 4.800 39.900 ;
        RECT 3.800 37.900 4.800 38.200 ;
        RECT 6.600 37.900 7.000 39.900 ;
        RECT 8.700 37.900 9.300 39.900 ;
        RECT 3.800 37.500 4.200 37.900 ;
        RECT 6.600 37.600 6.900 37.900 ;
        RECT 5.500 37.300 7.300 37.600 ;
        RECT 8.600 37.500 9.000 37.900 ;
        RECT 5.500 37.200 5.900 37.300 ;
        RECT 6.900 37.200 7.300 37.300 ;
        RECT 3.800 36.500 4.200 36.600 ;
        RECT 6.100 36.500 6.500 36.600 ;
        RECT 3.800 36.200 6.500 36.500 ;
        RECT 6.800 36.500 7.900 36.800 ;
        RECT 6.800 35.900 7.100 36.500 ;
        RECT 7.500 36.400 7.900 36.500 ;
        RECT 8.700 36.600 9.400 37.000 ;
        RECT 8.700 36.100 9.000 36.600 ;
        RECT 4.700 35.700 7.100 35.900 ;
        RECT 2.200 35.600 7.100 35.700 ;
        RECT 7.800 35.800 9.000 36.100 ;
        RECT 2.200 35.500 5.100 35.600 ;
        RECT 2.200 35.400 5.000 35.500 ;
        RECT 5.400 35.100 5.800 35.200 ;
        RECT 0.600 34.800 1.800 35.100 ;
        RECT 0.600 32.400 1.000 33.200 ;
        RECT 1.400 31.100 1.800 34.800 ;
        RECT 3.300 34.800 5.800 35.100 ;
        RECT 3.300 34.700 3.700 34.800 ;
        RECT 4.100 34.200 4.500 34.300 ;
        RECT 7.800 34.200 8.100 35.800 ;
        RECT 11.000 35.600 11.400 39.900 ;
        RECT 13.700 36.400 14.100 39.900 ;
        RECT 15.800 37.500 16.200 39.500 ;
        RECT 13.300 36.100 14.100 36.400 ;
        RECT 9.300 35.300 11.400 35.600 ;
        RECT 9.300 35.200 9.700 35.300 ;
        RECT 10.100 34.900 10.500 35.000 ;
        RECT 8.600 34.600 10.500 34.900 ;
        RECT 8.600 34.500 9.000 34.600 ;
        RECT 2.600 33.900 8.100 34.200 ;
        RECT 2.600 33.800 3.400 33.900 ;
        RECT 2.200 31.100 2.600 33.500 ;
        RECT 4.700 32.800 5.000 33.900 ;
        RECT 6.200 33.800 6.600 33.900 ;
        RECT 7.500 33.800 7.900 33.900 ;
        RECT 11.000 33.600 11.400 35.300 ;
        RECT 12.600 34.800 13.000 35.600 ;
        RECT 13.300 34.200 13.600 36.100 ;
        RECT 15.900 35.800 16.200 37.500 ;
        RECT 14.300 35.500 16.200 35.800 ;
        RECT 14.300 34.500 14.600 35.500 ;
        RECT 12.600 33.800 13.600 34.200 ;
        RECT 13.900 34.100 14.600 34.500 ;
        RECT 15.000 34.400 15.400 35.200 ;
        RECT 15.800 34.400 16.200 35.200 ;
        RECT 9.500 33.300 11.400 33.600 ;
        RECT 9.500 33.200 9.900 33.300 ;
        RECT 3.800 32.100 4.200 32.500 ;
        RECT 4.600 32.400 5.000 32.800 ;
        RECT 5.500 32.700 5.900 32.800 ;
        RECT 5.500 32.400 6.900 32.700 ;
        RECT 6.600 32.100 6.900 32.400 ;
        RECT 8.600 32.100 9.000 32.500 ;
        RECT 3.800 31.800 4.800 32.100 ;
        RECT 4.400 31.100 4.800 31.800 ;
        RECT 6.600 31.100 7.000 32.100 ;
        RECT 8.600 31.800 9.300 32.100 ;
        RECT 8.700 31.100 9.300 31.800 ;
        RECT 11.000 31.100 11.400 33.300 ;
        RECT 13.300 33.500 13.600 33.800 ;
        RECT 14.100 33.900 14.600 34.100 ;
        RECT 16.600 34.100 17.000 34.200 ;
        RECT 17.400 34.100 17.800 39.900 ;
        RECT 18.200 37.500 18.600 39.500 ;
        RECT 18.200 35.800 18.500 37.500 ;
        RECT 20.300 36.400 20.700 39.900 ;
        RECT 20.300 36.100 21.100 36.400 ;
        RECT 18.200 35.500 20.100 35.800 ;
        RECT 18.200 34.400 18.600 35.200 ;
        RECT 19.000 34.400 19.400 35.200 ;
        RECT 19.800 34.500 20.100 35.500 ;
        RECT 14.100 33.600 16.200 33.900 ;
        RECT 16.600 33.800 17.800 34.100 ;
        RECT 19.800 34.100 20.500 34.500 ;
        RECT 20.800 34.200 21.100 36.100 ;
        RECT 23.000 35.700 23.400 39.900 ;
        RECT 25.200 38.200 25.600 39.900 ;
        RECT 24.600 37.900 25.600 38.200 ;
        RECT 27.400 37.900 27.800 39.900 ;
        RECT 29.500 37.900 30.100 39.900 ;
        RECT 24.600 37.500 25.000 37.900 ;
        RECT 27.400 37.600 27.700 37.900 ;
        RECT 26.300 37.300 28.100 37.600 ;
        RECT 29.400 37.500 29.800 37.900 ;
        RECT 26.300 37.200 26.700 37.300 ;
        RECT 27.700 37.200 28.100 37.300 ;
        RECT 24.600 36.500 25.000 36.600 ;
        RECT 26.900 36.500 27.300 36.600 ;
        RECT 24.600 36.200 27.300 36.500 ;
        RECT 27.600 36.500 28.700 36.800 ;
        RECT 27.600 35.900 27.900 36.500 ;
        RECT 28.300 36.400 28.700 36.500 ;
        RECT 29.500 36.600 30.200 37.000 ;
        RECT 29.500 36.100 29.800 36.600 ;
        RECT 25.500 35.700 27.900 35.900 ;
        RECT 23.000 35.600 27.900 35.700 ;
        RECT 28.600 35.800 29.800 36.100 ;
        RECT 21.400 35.100 21.800 35.600 ;
        RECT 23.000 35.500 25.900 35.600 ;
        RECT 23.000 35.400 25.800 35.500 ;
        RECT 22.200 35.100 22.600 35.200 ;
        RECT 26.200 35.100 26.600 35.200 ;
        RECT 27.000 35.100 27.400 35.200 ;
        RECT 21.400 34.800 22.600 35.100 ;
        RECT 24.100 34.800 27.400 35.100 ;
        RECT 24.100 34.700 24.500 34.800 ;
        RECT 24.900 34.200 25.300 34.300 ;
        RECT 28.600 34.200 28.900 35.800 ;
        RECT 31.800 35.600 32.200 39.900 ;
        RECT 33.900 36.200 34.300 39.900 ;
        RECT 34.600 36.800 35.000 37.200 ;
        RECT 34.700 36.200 35.000 36.800 ;
        RECT 33.900 35.900 34.400 36.200 ;
        RECT 34.700 36.100 35.400 36.200 ;
        RECT 36.600 36.100 37.000 39.900 ;
        RECT 34.700 35.900 37.000 36.100 ;
        RECT 30.100 35.300 32.200 35.600 ;
        RECT 30.100 35.200 30.500 35.300 ;
        RECT 30.900 34.900 31.300 35.000 ;
        RECT 29.400 34.600 31.300 34.900 ;
        RECT 29.400 34.500 29.800 34.600 ;
        RECT 19.800 33.900 20.300 34.100 ;
        RECT 13.300 33.300 13.700 33.500 ;
        RECT 13.300 33.000 14.100 33.300 ;
        RECT 13.700 32.200 14.100 33.000 ;
        RECT 15.900 32.500 16.200 33.600 ;
        RECT 13.400 31.800 14.100 32.200 ;
        RECT 13.700 31.500 14.100 31.800 ;
        RECT 15.800 31.500 16.200 32.500 ;
        RECT 16.600 32.400 17.000 33.200 ;
        RECT 17.400 31.100 17.800 33.800 ;
        RECT 18.200 33.600 20.300 33.900 ;
        RECT 20.800 33.800 21.800 34.200 ;
        RECT 23.400 33.900 28.900 34.200 ;
        RECT 23.400 33.800 24.200 33.900 ;
        RECT 18.200 32.500 18.500 33.600 ;
        RECT 20.800 33.500 21.100 33.800 ;
        RECT 20.700 33.300 21.100 33.500 ;
        RECT 20.300 33.000 21.100 33.300 ;
        RECT 18.200 31.500 18.600 32.500 ;
        RECT 20.300 32.200 20.700 33.000 ;
        RECT 20.300 31.800 21.000 32.200 ;
        RECT 20.300 31.500 20.700 31.800 ;
        RECT 23.000 31.100 23.400 33.500 ;
        RECT 25.500 33.200 25.800 33.900 ;
        RECT 28.300 33.800 28.700 33.900 ;
        RECT 31.800 33.600 32.200 35.300 ;
        RECT 34.100 35.200 34.400 35.900 ;
        RECT 35.000 35.800 37.000 35.900 ;
        RECT 37.400 35.800 37.800 36.600 ;
        RECT 33.400 34.400 33.800 35.200 ;
        RECT 34.100 34.800 34.600 35.200 ;
        RECT 34.100 34.200 34.400 34.800 ;
        RECT 32.600 34.100 33.000 34.200 ;
        RECT 32.600 33.800 33.400 34.100 ;
        RECT 34.100 33.800 35.400 34.200 ;
        RECT 33.000 33.600 33.400 33.800 ;
        RECT 30.300 33.300 32.200 33.600 ;
        RECT 30.300 33.200 30.700 33.300 ;
        RECT 24.600 32.100 25.000 32.500 ;
        RECT 25.400 32.400 25.800 33.200 ;
        RECT 26.300 32.700 26.700 32.800 ;
        RECT 26.300 32.400 27.700 32.700 ;
        RECT 27.400 32.100 27.700 32.400 ;
        RECT 29.400 32.100 29.800 32.500 ;
        RECT 24.600 31.800 25.600 32.100 ;
        RECT 25.200 31.100 25.600 31.800 ;
        RECT 27.400 31.100 27.800 32.100 ;
        RECT 29.400 31.800 30.100 32.100 ;
        RECT 29.500 31.100 30.100 31.800 ;
        RECT 31.800 31.100 32.200 33.300 ;
        RECT 32.700 33.100 34.500 33.300 ;
        RECT 35.000 33.100 35.300 33.800 ;
        RECT 35.800 33.400 36.200 34.200 ;
        RECT 36.600 33.100 37.000 35.800 ;
        RECT 32.600 33.000 34.600 33.100 ;
        RECT 32.600 31.100 33.000 33.000 ;
        RECT 34.200 31.100 34.600 33.000 ;
        RECT 35.000 31.100 35.400 33.100 ;
        RECT 36.600 32.800 37.500 33.100 ;
        RECT 37.100 31.100 37.500 32.800 ;
        RECT 38.200 32.400 38.600 33.200 ;
        RECT 39.000 31.100 39.400 39.900 ;
        RECT 39.800 36.200 40.200 39.900 ;
        RECT 41.400 36.200 41.800 39.900 ;
        RECT 39.800 35.900 41.800 36.200 ;
        RECT 42.200 35.900 42.600 39.900 ;
        RECT 44.300 39.200 44.700 39.900 ;
        RECT 43.800 38.800 44.700 39.200 ;
        RECT 44.300 36.200 44.700 38.800 ;
        RECT 45.000 36.800 45.400 37.200 ;
        RECT 45.100 36.200 45.400 36.800 ;
        RECT 46.200 36.200 46.600 39.900 ;
        RECT 47.800 36.200 48.200 39.900 ;
        RECT 44.300 35.900 44.800 36.200 ;
        RECT 45.100 35.900 45.800 36.200 ;
        RECT 46.200 35.900 48.200 36.200 ;
        RECT 48.600 35.900 49.000 39.900 ;
        RECT 51.000 36.200 51.400 39.900 ;
        RECT 52.600 36.200 53.000 39.900 ;
        RECT 51.000 35.900 53.000 36.200 ;
        RECT 53.400 35.900 53.800 39.900 ;
        RECT 55.500 39.200 55.900 39.900 ;
        RECT 55.000 38.800 55.900 39.200 ;
        RECT 55.500 36.300 55.900 38.800 ;
        RECT 57.900 39.200 58.300 39.900 ;
        RECT 57.900 38.800 58.600 39.200 ;
        RECT 57.900 36.300 58.300 38.800 ;
        RECT 55.000 35.900 55.900 36.300 ;
        RECT 57.400 35.900 58.300 36.300 ;
        RECT 59.400 36.800 59.800 37.200 ;
        RECT 59.400 36.200 59.700 36.800 ;
        RECT 60.100 36.200 60.500 39.900 ;
        RECT 63.000 36.400 63.400 39.900 ;
        RECT 59.000 35.900 59.700 36.200 ;
        RECT 60.000 35.900 60.500 36.200 ;
        RECT 40.200 35.200 40.600 35.400 ;
        RECT 42.200 35.200 42.500 35.900 ;
        RECT 39.800 34.900 40.600 35.200 ;
        RECT 41.400 34.900 42.600 35.200 ;
        RECT 39.800 34.800 40.200 34.900 ;
        RECT 40.600 33.800 41.000 34.600 ;
        RECT 41.400 33.100 41.700 34.900 ;
        RECT 42.200 34.800 42.600 34.900 ;
        RECT 43.800 34.400 44.200 35.200 ;
        RECT 44.500 34.200 44.800 35.900 ;
        RECT 45.400 35.800 45.800 35.900 ;
        RECT 46.600 35.200 47.000 35.400 ;
        RECT 48.600 35.200 48.900 35.900 ;
        RECT 51.400 35.200 51.800 35.400 ;
        RECT 53.400 35.200 53.700 35.900 ;
        RECT 46.200 34.900 47.000 35.200 ;
        RECT 47.800 34.900 49.000 35.200 ;
        RECT 46.200 34.800 46.600 34.900 ;
        RECT 47.800 34.800 48.200 34.900 ;
        RECT 48.600 34.800 49.000 34.900 ;
        RECT 51.000 34.900 51.800 35.200 ;
        RECT 52.600 34.900 53.800 35.200 ;
        RECT 51.000 34.800 51.400 34.900 ;
        RECT 43.000 34.100 43.400 34.200 ;
        RECT 43.000 33.800 43.800 34.100 ;
        RECT 44.500 33.800 45.800 34.200 ;
        RECT 47.000 33.800 47.400 34.600 ;
        RECT 43.400 33.600 43.800 33.800 ;
        RECT 41.400 31.100 41.800 33.100 ;
        RECT 42.200 32.800 42.600 33.200 ;
        RECT 43.100 33.100 44.900 33.300 ;
        RECT 45.400 33.100 45.700 33.800 ;
        RECT 47.800 33.100 48.100 34.800 ;
        RECT 51.800 33.800 52.200 34.600 ;
        RECT 43.000 33.000 45.000 33.100 ;
        RECT 42.100 32.400 42.500 32.800 ;
        RECT 43.000 31.100 43.400 33.000 ;
        RECT 44.600 31.100 45.000 33.000 ;
        RECT 45.400 31.100 45.800 33.100 ;
        RECT 47.800 31.100 48.200 33.100 ;
        RECT 48.600 32.800 49.000 33.200 ;
        RECT 52.600 33.100 52.900 34.900 ;
        RECT 53.400 34.800 53.800 34.900 ;
        RECT 55.100 34.200 55.400 35.900 ;
        RECT 55.800 34.800 56.200 35.600 ;
        RECT 57.500 34.200 57.800 35.900 ;
        RECT 59.000 35.800 59.400 35.900 ;
        RECT 58.200 35.100 58.600 35.600 ;
        RECT 59.000 35.100 59.300 35.800 ;
        RECT 58.200 34.800 59.300 35.100 ;
        RECT 60.000 34.200 60.300 35.900 ;
        RECT 62.900 35.800 63.400 36.400 ;
        RECT 64.600 36.200 65.000 39.900 ;
        RECT 63.700 35.900 65.000 36.200 ;
        RECT 66.700 36.200 67.100 39.900 ;
        RECT 67.400 36.800 67.800 37.200 ;
        RECT 67.500 36.200 67.800 36.800 ;
        RECT 66.700 35.900 67.200 36.200 ;
        RECT 67.500 35.900 68.200 36.200 ;
        RECT 60.600 35.100 61.000 35.200 ;
        RECT 61.400 35.100 61.800 35.200 ;
        RECT 60.600 34.800 61.800 35.100 ;
        RECT 60.600 34.400 61.000 34.800 ;
        RECT 62.900 34.200 63.200 35.800 ;
        RECT 63.700 34.900 64.000 35.900 ;
        RECT 66.900 35.200 67.200 35.900 ;
        RECT 67.800 35.800 68.200 35.900 ;
        RECT 68.600 35.800 69.000 36.600 ;
        RECT 63.500 34.500 64.000 34.900 ;
        RECT 55.000 33.800 55.400 34.200 ;
        RECT 57.400 33.800 57.800 34.200 ;
        RECT 59.000 34.100 60.300 34.200 ;
        RECT 61.400 34.100 61.800 34.200 ;
        RECT 48.500 32.400 48.900 32.800 ;
        RECT 52.600 31.100 53.000 33.100 ;
        RECT 53.400 32.800 53.800 33.200 ;
        RECT 53.300 32.400 53.700 32.800 ;
        RECT 54.200 32.400 54.600 33.200 ;
        RECT 55.100 32.100 55.400 33.800 ;
        RECT 56.600 32.400 57.000 33.200 ;
        RECT 57.500 32.100 57.800 33.800 ;
        RECT 58.200 33.800 60.300 34.100 ;
        RECT 61.000 33.800 61.800 34.100 ;
        RECT 62.200 34.100 62.600 34.200 ;
        RECT 62.900 34.100 63.400 34.200 ;
        RECT 62.200 33.800 63.400 34.100 ;
        RECT 58.200 33.200 58.500 33.800 ;
        RECT 58.200 32.800 58.600 33.200 ;
        RECT 59.100 33.100 59.400 33.800 ;
        RECT 61.000 33.600 61.400 33.800 ;
        RECT 59.900 33.100 61.700 33.300 ;
        RECT 62.900 33.100 63.200 33.800 ;
        RECT 63.700 33.700 64.000 34.500 ;
        RECT 64.500 34.800 65.000 35.200 ;
        RECT 64.500 34.400 64.900 34.800 ;
        RECT 66.200 34.400 66.600 35.200 ;
        RECT 66.900 34.800 67.400 35.200 ;
        RECT 67.800 35.100 68.100 35.800 ;
        RECT 69.400 35.100 69.800 39.900 ;
        RECT 71.800 36.400 72.200 39.900 ;
        RECT 67.800 34.800 69.800 35.100 ;
        RECT 66.900 34.200 67.200 34.800 ;
        RECT 65.400 34.100 65.800 34.200 ;
        RECT 65.400 33.800 66.200 34.100 ;
        RECT 66.900 33.800 68.200 34.200 ;
        RECT 63.700 33.400 65.000 33.700 ;
        RECT 65.800 33.600 66.200 33.800 ;
        RECT 55.000 31.100 55.400 32.100 ;
        RECT 57.400 31.100 57.800 32.100 ;
        RECT 59.000 31.100 59.400 33.100 ;
        RECT 59.800 33.000 61.800 33.100 ;
        RECT 59.800 31.100 60.200 33.000 ;
        RECT 61.400 31.100 61.800 33.000 ;
        RECT 62.900 32.800 63.400 33.100 ;
        RECT 63.000 31.100 63.400 32.800 ;
        RECT 64.600 31.100 65.000 33.400 ;
        RECT 65.500 33.100 67.300 33.300 ;
        RECT 67.800 33.100 68.100 33.800 ;
        RECT 69.400 33.100 69.800 34.800 ;
        RECT 71.700 35.900 72.200 36.400 ;
        RECT 73.400 36.200 73.800 39.900 ;
        RECT 72.500 35.900 73.800 36.200 ;
        RECT 71.700 34.200 72.000 35.900 ;
        RECT 72.500 34.900 72.800 35.900 ;
        RECT 75.000 35.600 75.400 39.900 ;
        RECT 76.600 35.600 77.000 39.900 ;
        RECT 79.500 39.200 79.900 39.900 ;
        RECT 79.500 38.800 80.200 39.200 ;
        RECT 79.500 36.300 79.900 38.800 ;
        RECT 79.000 35.900 79.900 36.300 ;
        RECT 81.000 36.800 81.400 37.200 ;
        RECT 81.000 36.200 81.300 36.800 ;
        RECT 81.700 36.200 82.100 39.900 ;
        RECT 80.600 35.900 81.300 36.200 ;
        RECT 81.600 35.900 82.100 36.200 ;
        RECT 85.100 36.200 85.500 39.900 ;
        RECT 85.800 36.800 86.200 37.200 ;
        RECT 85.900 36.200 86.200 36.800 ;
        RECT 85.100 35.900 85.600 36.200 ;
        RECT 85.900 35.900 86.600 36.200 ;
        RECT 75.000 35.200 77.000 35.600 ;
        RECT 72.300 34.500 72.800 34.900 ;
        RECT 70.200 33.400 70.600 34.200 ;
        RECT 71.700 33.800 72.200 34.200 ;
        RECT 65.400 33.000 67.400 33.100 ;
        RECT 65.400 31.100 65.800 33.000 ;
        RECT 67.000 31.100 67.400 33.000 ;
        RECT 67.800 31.100 68.200 33.100 ;
        RECT 68.900 32.800 69.800 33.100 ;
        RECT 71.700 33.100 72.000 33.800 ;
        RECT 72.500 33.700 72.800 34.500 ;
        RECT 73.300 34.800 73.800 35.200 ;
        RECT 73.300 34.400 73.700 34.800 ;
        RECT 75.000 33.800 75.400 35.200 ;
        RECT 79.100 34.200 79.400 35.900 ;
        RECT 80.600 35.800 81.000 35.900 ;
        RECT 79.800 34.800 80.200 35.600 ;
        RECT 81.600 35.200 81.900 35.900 ;
        RECT 81.400 34.800 81.900 35.200 ;
        RECT 81.600 34.200 81.900 34.800 ;
        RECT 82.200 34.400 82.600 35.200 ;
        RECT 84.600 34.400 85.000 35.200 ;
        RECT 85.300 34.200 85.600 35.900 ;
        RECT 86.200 35.800 86.600 35.900 ;
        RECT 87.000 35.800 87.400 36.600 ;
        RECT 86.200 35.100 86.500 35.800 ;
        RECT 87.800 35.100 88.200 39.900 ;
        RECT 86.200 34.800 88.200 35.100 ;
        RECT 72.500 33.400 73.800 33.700 ;
        RECT 71.700 32.800 72.200 33.100 ;
        RECT 68.900 31.100 69.300 32.800 ;
        RECT 71.800 31.100 72.200 32.800 ;
        RECT 73.400 31.100 73.800 33.400 ;
        RECT 75.000 33.400 77.000 33.800 ;
        RECT 77.400 33.400 77.800 34.200 ;
        RECT 79.000 33.800 79.400 34.200 ;
        RECT 80.600 33.800 81.900 34.200 ;
        RECT 83.000 34.100 83.400 34.200 ;
        RECT 82.600 33.800 83.400 34.100 ;
        RECT 83.800 34.100 84.200 34.200 ;
        RECT 83.800 33.800 84.600 34.100 ;
        RECT 85.300 33.800 86.600 34.200 ;
        RECT 75.000 31.100 75.400 33.400 ;
        RECT 76.600 31.100 77.000 33.400 ;
        RECT 78.200 32.400 78.600 33.200 ;
        RECT 79.100 32.100 79.400 33.800 ;
        RECT 80.700 33.100 81.000 33.800 ;
        RECT 82.600 33.600 83.000 33.800 ;
        RECT 84.200 33.600 84.600 33.800 ;
        RECT 81.500 33.100 83.300 33.300 ;
        RECT 83.900 33.100 85.700 33.300 ;
        RECT 86.200 33.100 86.500 33.800 ;
        RECT 87.800 33.100 88.200 34.800 ;
        RECT 89.400 35.600 89.800 39.900 ;
        RECT 91.500 37.900 92.100 39.900 ;
        RECT 93.800 37.900 94.200 39.900 ;
        RECT 96.000 38.200 96.400 39.900 ;
        RECT 96.000 37.900 97.000 38.200 ;
        RECT 91.800 37.500 92.200 37.900 ;
        RECT 93.900 37.600 94.200 37.900 ;
        RECT 93.500 37.300 95.300 37.600 ;
        RECT 96.600 37.500 97.000 37.900 ;
        RECT 93.500 37.200 93.900 37.300 ;
        RECT 94.900 37.200 95.300 37.300 ;
        RECT 91.400 36.600 92.100 37.000 ;
        RECT 91.800 36.100 92.100 36.600 ;
        RECT 92.900 36.500 94.000 36.800 ;
        RECT 92.900 36.400 93.300 36.500 ;
        RECT 91.800 35.800 93.000 36.100 ;
        RECT 89.400 35.300 91.500 35.600 ;
        RECT 88.600 34.100 89.000 34.200 ;
        RECT 89.400 34.100 89.800 35.300 ;
        RECT 91.100 35.200 91.500 35.300 ;
        RECT 90.300 34.900 90.700 35.000 ;
        RECT 90.300 34.600 92.200 34.900 ;
        RECT 91.800 34.500 92.200 34.600 ;
        RECT 88.600 33.800 89.800 34.100 ;
        RECT 92.700 34.200 93.000 35.800 ;
        RECT 93.700 35.900 94.000 36.500 ;
        RECT 94.300 36.500 94.700 36.600 ;
        RECT 96.600 36.500 97.000 36.600 ;
        RECT 94.300 36.200 97.000 36.500 ;
        RECT 93.700 35.700 96.100 35.900 ;
        RECT 98.200 35.700 98.600 39.900 ;
        RECT 99.300 36.300 99.700 39.900 ;
        RECT 99.300 35.900 100.200 36.300 ;
        RECT 104.300 35.900 105.300 39.900 ;
        RECT 108.900 37.200 109.300 39.900 ;
        RECT 111.000 37.500 111.400 39.500 ;
        RECT 108.600 36.800 109.300 37.200 ;
        RECT 108.900 36.400 109.300 36.800 ;
        RECT 108.500 36.100 109.300 36.400 ;
        RECT 93.700 35.600 98.600 35.700 ;
        RECT 95.700 35.500 98.600 35.600 ;
        RECT 95.800 35.400 98.600 35.500 ;
        RECT 93.400 35.100 93.800 35.200 ;
        RECT 95.000 35.100 95.400 35.200 ;
        RECT 93.400 34.800 97.500 35.100 ;
        RECT 99.000 34.800 99.400 35.600 ;
        RECT 97.100 34.700 97.500 34.800 ;
        RECT 96.300 34.200 96.700 34.300 ;
        RECT 99.800 34.200 100.100 35.900 ;
        RECT 103.800 34.400 104.200 35.200 ;
        RECT 104.600 34.200 104.900 35.900 ;
        RECT 105.400 34.400 105.800 35.200 ;
        RECT 107.800 34.800 108.200 35.600 ;
        RECT 92.700 33.900 98.200 34.200 ;
        RECT 92.900 33.800 93.300 33.900 ;
        RECT 88.600 33.400 89.000 33.800 ;
        RECT 89.400 33.600 89.800 33.800 ;
        RECT 79.000 31.100 79.400 32.100 ;
        RECT 80.600 31.100 81.000 33.100 ;
        RECT 81.400 33.000 83.400 33.100 ;
        RECT 81.400 31.100 81.800 33.000 ;
        RECT 83.000 31.100 83.400 33.000 ;
        RECT 83.800 33.000 85.800 33.100 ;
        RECT 83.800 31.100 84.200 33.000 ;
        RECT 85.400 31.100 85.800 33.000 ;
        RECT 86.200 31.100 86.600 33.100 ;
        RECT 87.300 32.800 88.200 33.100 ;
        RECT 89.400 33.300 91.300 33.600 ;
        RECT 87.300 31.100 87.700 32.800 ;
        RECT 89.400 31.100 89.800 33.300 ;
        RECT 90.900 33.200 91.300 33.300 ;
        RECT 95.800 32.800 96.100 33.900 ;
        RECT 97.400 33.800 98.200 33.900 ;
        RECT 99.800 34.100 100.200 34.200 ;
        RECT 103.000 34.100 103.400 34.200 ;
        RECT 104.600 34.100 105.000 34.200 ;
        RECT 99.800 33.800 103.800 34.100 ;
        RECT 104.600 33.800 105.800 34.100 ;
        RECT 106.200 33.800 106.600 34.600 ;
        RECT 108.500 34.200 108.800 36.100 ;
        RECT 111.100 35.800 111.400 37.500 ;
        RECT 111.800 36.200 112.200 39.900 ;
        RECT 113.400 36.200 113.800 39.900 ;
        RECT 111.800 35.900 113.800 36.200 ;
        RECT 114.200 35.900 114.600 39.900 ;
        RECT 109.500 35.500 111.400 35.800 ;
        RECT 109.500 34.500 109.800 35.500 ;
        RECT 112.200 35.200 112.600 35.400 ;
        RECT 114.200 35.200 114.500 35.900 ;
        RECT 107.800 33.800 108.800 34.200 ;
        RECT 109.100 34.100 109.800 34.500 ;
        RECT 110.200 34.400 110.600 35.200 ;
        RECT 111.000 34.400 111.400 35.200 ;
        RECT 111.800 34.900 112.600 35.200 ;
        RECT 113.400 34.900 114.600 35.200 ;
        RECT 111.800 34.800 112.200 34.900 ;
        RECT 94.900 32.700 95.300 32.800 ;
        RECT 91.800 32.100 92.200 32.500 ;
        RECT 93.900 32.400 95.300 32.700 ;
        RECT 95.800 32.400 96.200 32.800 ;
        RECT 93.900 32.100 94.200 32.400 ;
        RECT 96.600 32.100 97.000 32.500 ;
        RECT 91.500 31.800 92.200 32.100 ;
        RECT 91.500 31.100 92.100 31.800 ;
        RECT 93.800 31.100 94.200 32.100 ;
        RECT 96.000 31.800 97.000 32.100 ;
        RECT 96.000 31.100 96.400 31.800 ;
        RECT 98.200 31.100 98.600 33.500 ;
        RECT 99.800 32.100 100.100 33.800 ;
        RECT 103.400 33.600 103.800 33.800 ;
        RECT 100.600 32.400 101.000 33.200 ;
        RECT 103.100 33.100 104.900 33.300 ;
        RECT 105.500 33.100 105.800 33.800 ;
        RECT 108.500 33.500 108.800 33.800 ;
        RECT 109.300 33.900 109.800 34.100 ;
        RECT 109.300 33.600 111.400 33.900 ;
        RECT 112.600 33.800 113.000 34.600 ;
        RECT 108.500 33.300 108.900 33.500 ;
        RECT 103.000 33.000 105.000 33.100 ;
        RECT 99.800 31.100 100.200 32.100 ;
        RECT 103.000 31.100 103.400 33.000 ;
        RECT 104.600 31.400 105.000 33.000 ;
        RECT 105.400 31.700 105.800 33.100 ;
        RECT 106.200 31.400 106.600 33.100 ;
        RECT 108.500 33.000 109.300 33.300 ;
        RECT 108.900 31.500 109.300 33.000 ;
        RECT 111.100 32.500 111.400 33.600 ;
        RECT 111.000 31.500 111.400 32.500 ;
        RECT 113.400 33.100 113.700 34.900 ;
        RECT 114.200 34.800 114.600 34.900 ;
        RECT 115.000 34.100 115.400 39.900 ;
        RECT 116.600 35.600 117.000 39.900 ;
        RECT 118.700 37.900 119.300 39.900 ;
        RECT 121.000 37.900 121.400 39.900 ;
        RECT 123.200 38.200 123.600 39.900 ;
        RECT 123.200 37.900 124.200 38.200 ;
        RECT 119.000 37.500 119.400 37.900 ;
        RECT 121.100 37.600 121.400 37.900 ;
        RECT 120.700 37.300 122.500 37.600 ;
        RECT 123.800 37.500 124.200 37.900 ;
        RECT 120.700 37.200 121.100 37.300 ;
        RECT 122.100 37.200 122.500 37.300 ;
        RECT 118.600 36.600 119.300 37.000 ;
        RECT 119.000 36.100 119.300 36.600 ;
        RECT 120.100 36.500 121.200 36.800 ;
        RECT 120.100 36.400 120.500 36.500 ;
        RECT 119.000 35.800 120.200 36.100 ;
        RECT 116.600 35.300 118.700 35.600 ;
        RECT 115.800 34.100 116.200 34.200 ;
        RECT 115.000 33.800 116.200 34.100 ;
        RECT 104.600 31.100 106.600 31.400 ;
        RECT 113.400 31.100 113.800 33.100 ;
        RECT 114.200 32.800 114.600 33.200 ;
        RECT 114.100 32.400 114.500 32.800 ;
        RECT 115.000 31.100 115.400 33.800 ;
        RECT 116.600 33.600 117.000 35.300 ;
        RECT 118.300 35.200 118.700 35.300 ;
        RECT 117.500 34.900 117.900 35.000 ;
        RECT 117.500 34.600 119.400 34.900 ;
        RECT 119.000 34.500 119.400 34.600 ;
        RECT 119.900 34.200 120.200 35.800 ;
        RECT 120.900 35.900 121.200 36.500 ;
        RECT 121.500 36.500 121.900 36.600 ;
        RECT 123.800 36.500 124.200 36.600 ;
        RECT 121.500 36.200 124.200 36.500 ;
        RECT 120.900 35.700 123.300 35.900 ;
        RECT 125.400 35.700 125.800 39.900 ;
        RECT 127.500 36.300 127.900 39.900 ;
        RECT 127.000 35.900 127.900 36.300 ;
        RECT 128.600 35.900 129.000 39.900 ;
        RECT 129.400 36.200 129.800 39.900 ;
        RECT 131.000 36.200 131.400 39.900 ;
        RECT 133.700 36.400 134.100 39.900 ;
        RECT 135.800 37.500 136.200 39.500 ;
        RECT 129.400 35.900 131.400 36.200 ;
        RECT 133.300 36.100 134.100 36.400 ;
        RECT 120.900 35.600 125.800 35.700 ;
        RECT 122.900 35.500 125.800 35.600 ;
        RECT 123.000 35.400 125.800 35.500 ;
        RECT 120.600 35.100 121.000 35.200 ;
        RECT 122.200 35.100 122.600 35.200 ;
        RECT 120.600 34.800 124.700 35.100 ;
        RECT 124.300 34.700 124.700 34.800 ;
        RECT 123.500 34.200 123.900 34.300 ;
        RECT 127.100 34.200 127.400 35.900 ;
        RECT 127.800 34.800 128.200 35.600 ;
        RECT 128.700 35.200 129.000 35.900 ;
        RECT 130.600 35.200 131.000 35.400 ;
        RECT 128.600 34.900 129.800 35.200 ;
        RECT 130.600 35.100 131.400 35.200 ;
        RECT 132.600 35.100 133.000 35.600 ;
        RECT 130.600 34.900 133.000 35.100 ;
        RECT 128.600 34.800 129.000 34.900 ;
        RECT 119.900 33.900 125.400 34.200 ;
        RECT 120.100 33.800 120.500 33.900 ;
        RECT 116.600 33.300 118.500 33.600 ;
        RECT 115.800 33.100 116.200 33.200 ;
        RECT 116.600 33.100 117.000 33.300 ;
        RECT 118.100 33.200 118.500 33.300 ;
        RECT 115.800 32.800 117.000 33.100 ;
        RECT 123.000 32.800 123.300 33.900 ;
        RECT 124.600 33.800 125.400 33.900 ;
        RECT 127.000 33.800 127.400 34.200 ;
        RECT 115.800 32.400 116.200 32.800 ;
        RECT 116.600 31.100 117.000 32.800 ;
        RECT 122.100 32.700 122.500 32.800 ;
        RECT 119.000 32.100 119.400 32.500 ;
        RECT 121.100 32.400 122.500 32.700 ;
        RECT 123.000 32.400 123.400 32.800 ;
        RECT 121.100 32.100 121.400 32.400 ;
        RECT 123.800 32.100 124.200 32.500 ;
        RECT 118.700 31.800 119.400 32.100 ;
        RECT 118.700 31.100 119.300 31.800 ;
        RECT 121.000 31.100 121.400 32.100 ;
        RECT 123.200 31.800 124.200 32.100 ;
        RECT 123.200 31.100 123.600 31.800 ;
        RECT 125.400 31.100 125.800 33.500 ;
        RECT 126.200 32.400 126.600 33.200 ;
        RECT 127.100 33.100 127.400 33.800 ;
        RECT 128.600 33.100 129.000 33.200 ;
        RECT 129.500 33.100 129.800 34.900 ;
        RECT 131.000 34.800 133.000 34.900 ;
        RECT 133.300 35.200 133.600 36.100 ;
        RECT 135.900 35.800 136.200 37.500 ;
        RECT 134.300 35.500 136.200 35.800 ;
        RECT 136.600 37.100 137.000 39.900 ;
        RECT 137.400 37.100 137.800 37.200 ;
        RECT 136.600 36.800 137.800 37.100 ;
        RECT 133.300 34.800 133.800 35.200 ;
        RECT 130.200 33.800 130.600 34.600 ;
        RECT 133.300 34.200 133.600 34.800 ;
        RECT 134.300 34.500 134.600 35.500 ;
        RECT 132.600 33.800 133.600 34.200 ;
        RECT 133.900 34.100 134.600 34.500 ;
        RECT 135.000 34.400 135.400 35.200 ;
        RECT 135.800 34.400 136.200 35.200 ;
        RECT 127.000 32.800 129.000 33.100 ;
        RECT 127.100 32.100 127.400 32.800 ;
        RECT 128.700 32.400 129.100 32.800 ;
        RECT 127.000 31.100 127.400 32.100 ;
        RECT 129.400 31.100 129.800 33.100 ;
        RECT 133.300 33.500 133.600 33.800 ;
        RECT 134.100 33.900 134.600 34.100 ;
        RECT 134.100 33.600 136.200 33.900 ;
        RECT 133.300 33.300 133.700 33.500 ;
        RECT 133.300 33.000 134.100 33.300 ;
        RECT 133.700 31.500 134.100 33.000 ;
        RECT 135.900 32.500 136.200 33.600 ;
        RECT 135.800 31.500 136.200 32.500 ;
        RECT 136.600 31.100 137.000 36.800 ;
        RECT 138.200 35.600 138.600 39.900 ;
        RECT 140.300 37.900 140.900 39.900 ;
        RECT 142.600 37.900 143.000 39.900 ;
        RECT 144.800 38.200 145.200 39.900 ;
        RECT 144.800 37.900 145.800 38.200 ;
        RECT 140.600 37.500 141.000 37.900 ;
        RECT 142.700 37.600 143.000 37.900 ;
        RECT 142.300 37.300 144.100 37.600 ;
        RECT 145.400 37.500 145.800 37.900 ;
        RECT 142.300 37.200 142.700 37.300 ;
        RECT 143.700 37.200 144.100 37.300 ;
        RECT 139.800 37.000 140.500 37.200 ;
        RECT 139.800 36.800 140.900 37.000 ;
        RECT 140.200 36.600 140.900 36.800 ;
        RECT 140.600 36.100 140.900 36.600 ;
        RECT 141.700 36.500 142.800 36.800 ;
        RECT 141.700 36.400 142.100 36.500 ;
        RECT 140.600 35.800 141.800 36.100 ;
        RECT 138.200 35.300 140.300 35.600 ;
        RECT 138.200 33.600 138.600 35.300 ;
        RECT 139.900 35.200 140.300 35.300 ;
        RECT 139.100 34.900 139.500 35.000 ;
        RECT 139.100 34.600 141.000 34.900 ;
        RECT 140.600 34.500 141.000 34.600 ;
        RECT 141.500 34.200 141.800 35.800 ;
        RECT 142.500 35.900 142.800 36.500 ;
        RECT 143.100 36.500 143.500 36.600 ;
        RECT 145.400 36.500 145.800 36.600 ;
        RECT 143.100 36.200 145.800 36.500 ;
        RECT 142.500 35.700 144.900 35.900 ;
        RECT 147.000 35.700 147.400 39.900 ;
        RECT 142.500 35.600 147.400 35.700 ;
        RECT 148.600 35.600 149.000 39.900 ;
        RECT 150.200 35.600 150.600 39.900 ;
        RECT 151.800 35.600 152.200 39.900 ;
        RECT 153.400 35.600 153.800 39.900 ;
        RECT 144.500 35.500 147.400 35.600 ;
        RECT 144.600 35.400 147.400 35.500 ;
        RECT 147.800 35.200 149.000 35.600 ;
        RECT 149.500 35.200 150.600 35.600 ;
        RECT 151.100 35.200 152.200 35.600 ;
        RECT 152.900 35.200 153.800 35.600 ;
        RECT 142.200 35.100 142.600 35.200 ;
        RECT 143.800 35.100 144.200 35.200 ;
        RECT 142.200 34.800 146.300 35.100 ;
        RECT 145.900 34.700 146.300 34.800 ;
        RECT 145.100 34.200 145.500 34.300 ;
        RECT 141.500 33.900 147.000 34.200 ;
        RECT 141.700 33.800 142.100 33.900 ;
        RECT 138.200 33.300 140.100 33.600 ;
        RECT 137.400 33.100 137.800 33.200 ;
        RECT 138.200 33.100 138.600 33.300 ;
        RECT 139.700 33.200 140.100 33.300 ;
        RECT 137.400 32.800 138.600 33.100 ;
        RECT 144.600 32.800 144.900 33.900 ;
        RECT 146.200 33.800 147.000 33.900 ;
        RECT 147.800 33.800 148.200 35.200 ;
        RECT 149.500 34.500 149.900 35.200 ;
        RECT 151.100 34.500 151.500 35.200 ;
        RECT 152.900 34.500 153.300 35.200 ;
        RECT 148.600 34.100 149.900 34.500 ;
        RECT 150.300 34.100 151.500 34.500 ;
        RECT 152.000 34.100 153.300 34.500 ;
        RECT 149.500 33.800 149.900 34.100 ;
        RECT 151.100 33.800 151.500 34.100 ;
        RECT 152.900 33.800 153.300 34.100 ;
        RECT 137.400 32.400 137.800 32.800 ;
        RECT 138.200 31.100 138.600 32.800 ;
        RECT 143.700 32.700 144.100 32.800 ;
        RECT 140.600 32.100 141.000 32.500 ;
        RECT 142.700 32.400 144.100 32.700 ;
        RECT 144.600 32.400 145.000 32.800 ;
        RECT 142.700 32.100 143.000 32.400 ;
        RECT 145.400 32.100 145.800 32.500 ;
        RECT 140.300 31.800 141.000 32.100 ;
        RECT 140.300 31.100 140.900 31.800 ;
        RECT 142.600 31.100 143.000 32.100 ;
        RECT 144.800 31.800 145.800 32.100 ;
        RECT 144.800 31.100 145.200 31.800 ;
        RECT 147.000 31.100 147.400 33.500 ;
        RECT 147.800 33.400 149.000 33.800 ;
        RECT 149.500 33.400 150.600 33.800 ;
        RECT 151.100 33.400 152.200 33.800 ;
        RECT 152.900 33.400 153.800 33.800 ;
        RECT 148.600 31.100 149.000 33.400 ;
        RECT 150.200 31.100 150.600 33.400 ;
        RECT 151.800 31.100 152.200 33.400 ;
        RECT 153.400 31.100 153.800 33.400 ;
        RECT 156.600 31.100 157.000 39.900 ;
        RECT 158.200 35.600 158.600 39.900 ;
        RECT 160.300 37.900 160.900 39.900 ;
        RECT 162.600 37.900 163.000 39.900 ;
        RECT 164.800 38.200 165.200 39.900 ;
        RECT 164.800 37.900 165.800 38.200 ;
        RECT 160.600 37.500 161.000 37.900 ;
        RECT 162.700 37.600 163.000 37.900 ;
        RECT 162.300 37.300 164.100 37.600 ;
        RECT 165.400 37.500 165.800 37.900 ;
        RECT 162.300 37.200 162.700 37.300 ;
        RECT 163.700 37.200 164.100 37.300 ;
        RECT 160.200 36.600 160.900 37.000 ;
        RECT 160.600 36.100 160.900 36.600 ;
        RECT 161.700 36.500 162.800 36.800 ;
        RECT 161.700 36.400 162.100 36.500 ;
        RECT 160.600 35.800 161.800 36.100 ;
        RECT 158.200 35.300 160.300 35.600 ;
        RECT 158.200 33.600 158.600 35.300 ;
        RECT 159.900 35.200 160.300 35.300 ;
        RECT 159.100 34.900 159.500 35.000 ;
        RECT 159.100 34.600 161.000 34.900 ;
        RECT 160.600 34.500 161.000 34.600 ;
        RECT 161.500 34.200 161.800 35.800 ;
        RECT 162.500 35.900 162.800 36.500 ;
        RECT 163.100 36.500 163.500 36.600 ;
        RECT 165.400 36.500 165.800 36.600 ;
        RECT 163.100 36.200 165.800 36.500 ;
        RECT 162.500 35.700 164.900 35.900 ;
        RECT 167.000 35.700 167.400 39.900 ;
        RECT 169.100 36.300 169.500 39.900 ;
        RECT 168.600 35.900 169.500 36.300 ;
        RECT 170.200 35.900 170.600 39.900 ;
        RECT 171.000 36.200 171.400 39.900 ;
        RECT 172.600 36.200 173.000 39.900 ;
        RECT 171.000 35.900 173.000 36.200 ;
        RECT 173.400 37.500 173.800 39.500 ;
        RECT 162.500 35.600 167.400 35.700 ;
        RECT 164.500 35.500 167.400 35.600 ;
        RECT 164.600 35.400 167.400 35.500 ;
        RECT 162.200 35.100 162.600 35.200 ;
        RECT 163.800 35.100 164.200 35.200 ;
        RECT 162.200 34.800 166.300 35.100 ;
        RECT 165.900 34.700 166.300 34.800 ;
        RECT 165.100 34.200 165.500 34.300 ;
        RECT 168.700 34.200 169.000 35.900 ;
        RECT 169.400 34.800 169.800 35.600 ;
        RECT 170.300 35.200 170.600 35.900 ;
        RECT 173.400 35.800 173.700 37.500 ;
        RECT 175.500 36.400 175.900 39.900 ;
        RECT 175.500 36.100 176.300 36.400 ;
        RECT 173.400 35.500 175.300 35.800 ;
        RECT 172.200 35.200 172.600 35.400 ;
        RECT 170.200 34.900 171.400 35.200 ;
        RECT 172.200 34.900 173.000 35.200 ;
        RECT 170.200 34.800 170.600 34.900 ;
        RECT 161.500 33.900 167.000 34.200 ;
        RECT 161.700 33.800 162.100 33.900 ;
        RECT 158.200 33.300 160.100 33.600 ;
        RECT 157.400 33.100 157.800 33.200 ;
        RECT 158.200 33.100 158.600 33.300 ;
        RECT 159.700 33.200 160.100 33.300 ;
        RECT 157.400 32.800 158.600 33.100 ;
        RECT 164.600 32.800 164.900 33.900 ;
        RECT 166.200 33.800 167.000 33.900 ;
        RECT 168.600 33.800 169.000 34.200 ;
        RECT 157.400 32.400 157.800 32.800 ;
        RECT 158.200 31.100 158.600 32.800 ;
        RECT 163.700 32.700 164.100 32.800 ;
        RECT 160.600 32.100 161.000 32.500 ;
        RECT 162.700 32.400 164.100 32.700 ;
        RECT 164.600 32.400 165.000 32.800 ;
        RECT 162.700 32.100 163.000 32.400 ;
        RECT 165.400 32.100 165.800 32.500 ;
        RECT 160.300 31.800 161.000 32.100 ;
        RECT 160.300 31.100 160.900 31.800 ;
        RECT 162.600 31.100 163.000 32.100 ;
        RECT 164.800 31.800 165.800 32.100 ;
        RECT 164.800 31.100 165.200 31.800 ;
        RECT 167.000 31.100 167.400 33.500 ;
        RECT 167.800 32.400 168.200 33.200 ;
        RECT 168.700 33.100 169.000 33.800 ;
        RECT 170.200 33.100 170.600 33.200 ;
        RECT 171.100 33.100 171.400 34.900 ;
        RECT 172.600 34.800 173.000 34.900 ;
        RECT 171.800 33.800 172.200 34.600 ;
        RECT 173.400 34.400 173.800 35.200 ;
        RECT 174.200 34.400 174.600 35.200 ;
        RECT 175.000 34.500 175.300 35.500 ;
        RECT 175.000 34.100 175.700 34.500 ;
        RECT 176.000 34.200 176.300 36.100 ;
        RECT 178.200 36.100 178.600 39.900 ;
        RECT 181.100 36.300 181.500 39.900 ;
        RECT 179.000 36.100 179.400 36.200 ;
        RECT 178.200 35.800 179.400 36.100 ;
        RECT 180.600 35.900 181.500 36.300 ;
        RECT 182.200 35.900 182.600 39.900 ;
        RECT 183.000 36.200 183.400 39.900 ;
        RECT 184.600 36.200 185.000 39.900 ;
        RECT 183.000 35.900 185.000 36.200 ;
        RECT 176.600 34.800 177.000 35.600 ;
        RECT 176.000 34.100 177.000 34.200 ;
        RECT 177.400 34.100 177.800 34.200 ;
        RECT 175.000 33.900 175.500 34.100 ;
        RECT 168.600 32.800 170.600 33.100 ;
        RECT 168.700 32.100 169.000 32.800 ;
        RECT 170.300 32.400 170.700 32.800 ;
        RECT 168.600 31.100 169.000 32.100 ;
        RECT 171.000 31.100 171.400 33.100 ;
        RECT 173.400 33.600 175.500 33.900 ;
        RECT 176.000 33.800 177.800 34.100 ;
        RECT 173.400 32.500 173.700 33.600 ;
        RECT 176.000 33.500 176.300 33.800 ;
        RECT 175.900 33.300 176.300 33.500 ;
        RECT 175.500 33.000 176.300 33.300 ;
        RECT 173.400 31.500 173.800 32.500 ;
        RECT 175.500 31.500 175.900 33.000 ;
        RECT 178.200 31.100 178.600 35.800 ;
        RECT 180.700 34.200 181.000 35.900 ;
        RECT 181.400 34.800 181.800 35.600 ;
        RECT 182.300 35.200 182.600 35.900 ;
        RECT 185.400 35.600 185.800 39.900 ;
        RECT 187.500 37.900 188.100 39.900 ;
        RECT 189.800 37.900 190.200 39.900 ;
        RECT 192.000 38.200 192.400 39.900 ;
        RECT 192.000 37.900 193.000 38.200 ;
        RECT 187.800 37.500 188.200 37.900 ;
        RECT 189.900 37.600 190.200 37.900 ;
        RECT 189.500 37.300 191.300 37.600 ;
        RECT 192.600 37.500 193.000 37.900 ;
        RECT 189.500 37.200 189.900 37.300 ;
        RECT 190.900 37.200 191.300 37.300 ;
        RECT 187.400 36.600 188.100 37.000 ;
        RECT 187.800 36.100 188.100 36.600 ;
        RECT 188.900 36.500 190.000 36.800 ;
        RECT 188.900 36.400 189.300 36.500 ;
        RECT 187.800 35.800 189.000 36.100 ;
        RECT 184.200 35.200 184.600 35.400 ;
        RECT 185.400 35.300 187.500 35.600 ;
        RECT 182.200 34.900 183.400 35.200 ;
        RECT 184.200 34.900 185.000 35.200 ;
        RECT 182.200 34.800 182.600 34.900 ;
        RECT 180.600 33.800 181.000 34.200 ;
        RECT 179.000 32.400 179.400 33.200 ;
        RECT 179.800 32.400 180.200 33.200 ;
        RECT 180.700 33.100 181.000 33.800 ;
        RECT 182.200 33.100 182.600 33.200 ;
        RECT 183.100 33.100 183.400 34.900 ;
        RECT 184.600 34.800 185.000 34.900 ;
        RECT 183.800 33.800 184.200 34.600 ;
        RECT 184.600 34.100 185.000 34.200 ;
        RECT 185.400 34.100 185.800 35.300 ;
        RECT 187.100 35.200 187.500 35.300 ;
        RECT 188.700 35.200 189.000 35.800 ;
        RECT 189.700 35.900 190.000 36.500 ;
        RECT 190.300 36.500 190.700 36.600 ;
        RECT 192.600 36.500 193.000 36.600 ;
        RECT 190.300 36.200 193.000 36.500 ;
        RECT 189.700 35.700 192.100 35.900 ;
        RECT 194.200 35.700 194.600 39.900 ;
        RECT 189.700 35.600 194.600 35.700 ;
        RECT 191.700 35.500 194.600 35.600 ;
        RECT 191.800 35.400 194.600 35.500 ;
        RECT 195.000 35.600 195.400 39.900 ;
        RECT 197.100 37.900 197.700 39.900 ;
        RECT 199.400 37.900 199.800 39.900 ;
        RECT 201.600 38.200 202.000 39.900 ;
        RECT 201.600 37.900 202.600 38.200 ;
        RECT 197.400 37.500 197.800 37.900 ;
        RECT 199.500 37.600 199.800 37.900 ;
        RECT 199.100 37.300 200.900 37.600 ;
        RECT 202.200 37.500 202.600 37.900 ;
        RECT 199.100 37.200 199.500 37.300 ;
        RECT 200.500 37.200 200.900 37.300 ;
        RECT 197.000 36.600 197.700 37.000 ;
        RECT 197.400 36.100 197.700 36.600 ;
        RECT 198.500 36.500 199.600 36.800 ;
        RECT 198.500 36.400 198.900 36.500 ;
        RECT 197.400 35.800 198.600 36.100 ;
        RECT 195.000 35.300 197.100 35.600 ;
        RECT 186.300 34.900 186.700 35.000 ;
        RECT 186.300 34.600 188.200 34.900 ;
        RECT 188.600 34.800 189.000 35.200 ;
        RECT 189.400 35.100 189.800 35.200 ;
        RECT 191.000 35.100 191.400 35.200 ;
        RECT 189.400 34.800 193.500 35.100 ;
        RECT 187.800 34.500 188.200 34.600 ;
        RECT 184.600 33.800 185.800 34.100 ;
        RECT 188.700 34.200 189.000 34.800 ;
        RECT 193.100 34.700 193.500 34.800 ;
        RECT 192.300 34.200 192.700 34.300 ;
        RECT 188.700 33.900 194.200 34.200 ;
        RECT 188.900 33.800 189.300 33.900 ;
        RECT 180.600 32.800 182.600 33.100 ;
        RECT 180.700 32.100 181.000 32.800 ;
        RECT 182.300 32.400 182.700 32.800 ;
        RECT 180.600 31.100 181.000 32.100 ;
        RECT 183.000 31.100 183.400 33.100 ;
        RECT 185.400 33.600 185.800 33.800 ;
        RECT 185.400 33.300 187.300 33.600 ;
        RECT 185.400 31.100 185.800 33.300 ;
        RECT 186.900 33.200 187.300 33.300 ;
        RECT 191.800 32.800 192.100 33.900 ;
        RECT 193.400 33.800 194.200 33.900 ;
        RECT 195.000 33.600 195.400 35.300 ;
        RECT 196.700 35.200 197.100 35.300 ;
        RECT 198.300 35.200 198.600 35.800 ;
        RECT 199.300 35.900 199.600 36.500 ;
        RECT 199.900 36.500 200.300 36.600 ;
        RECT 202.200 36.500 202.600 36.600 ;
        RECT 199.900 36.200 202.600 36.500 ;
        RECT 199.300 35.700 201.700 35.900 ;
        RECT 203.800 35.700 204.200 39.900 ;
        RECT 199.300 35.600 204.200 35.700 ;
        RECT 201.300 35.500 204.200 35.600 ;
        RECT 201.400 35.400 204.200 35.500 ;
        RECT 195.900 34.900 196.300 35.000 ;
        RECT 195.900 34.600 197.800 34.900 ;
        RECT 198.200 34.800 198.600 35.200 ;
        RECT 200.600 35.100 201.000 35.200 ;
        RECT 200.600 34.800 203.100 35.100 ;
        RECT 197.400 34.500 197.800 34.600 ;
        RECT 198.300 34.200 198.600 34.800 ;
        RECT 201.400 34.700 201.800 34.800 ;
        RECT 202.700 34.700 203.100 34.800 ;
        RECT 201.900 34.200 202.300 34.300 ;
        RECT 198.300 33.900 203.800 34.200 ;
        RECT 198.500 33.800 198.900 33.900 ;
        RECT 190.900 32.700 191.300 32.800 ;
        RECT 187.800 32.100 188.200 32.500 ;
        RECT 189.900 32.400 191.300 32.700 ;
        RECT 191.800 32.400 192.200 32.800 ;
        RECT 189.900 32.100 190.200 32.400 ;
        RECT 192.600 32.100 193.000 32.500 ;
        RECT 187.500 31.800 188.200 32.100 ;
        RECT 187.500 31.100 188.100 31.800 ;
        RECT 189.800 31.100 190.200 32.100 ;
        RECT 192.000 31.800 193.000 32.100 ;
        RECT 192.000 31.100 192.400 31.800 ;
        RECT 194.200 31.100 194.600 33.500 ;
        RECT 195.000 33.300 196.900 33.600 ;
        RECT 195.000 31.100 195.400 33.300 ;
        RECT 196.500 33.200 196.900 33.300 ;
        RECT 201.400 32.800 201.700 33.900 ;
        RECT 203.000 33.800 203.800 33.900 ;
        RECT 200.500 32.700 200.900 32.800 ;
        RECT 197.400 32.100 197.800 32.500 ;
        RECT 199.500 32.400 200.900 32.700 ;
        RECT 201.400 32.400 201.800 32.800 ;
        RECT 199.500 32.100 199.800 32.400 ;
        RECT 202.200 32.100 202.600 32.500 ;
        RECT 197.100 31.800 197.800 32.100 ;
        RECT 197.100 31.100 197.700 31.800 ;
        RECT 199.400 31.100 199.800 32.100 ;
        RECT 201.600 31.800 202.600 32.100 ;
        RECT 201.600 31.100 202.000 31.800 ;
        RECT 203.800 31.100 204.200 33.500 ;
        RECT 0.600 27.700 1.000 29.900 ;
        RECT 2.700 29.200 3.300 29.900 ;
        RECT 2.700 28.900 3.400 29.200 ;
        RECT 5.000 28.900 5.400 29.900 ;
        RECT 7.200 29.200 7.600 29.900 ;
        RECT 7.200 28.900 8.200 29.200 ;
        RECT 3.000 28.500 3.400 28.900 ;
        RECT 5.100 28.600 5.400 28.900 ;
        RECT 5.100 28.300 6.500 28.600 ;
        RECT 6.100 28.200 6.500 28.300 ;
        RECT 7.000 28.200 7.400 28.600 ;
        RECT 7.800 28.500 8.200 28.900 ;
        RECT 2.100 27.700 2.500 27.800 ;
        RECT 0.600 27.400 2.500 27.700 ;
        RECT 0.600 25.700 1.000 27.400 ;
        RECT 4.100 27.100 4.500 27.200 ;
        RECT 6.200 27.100 6.600 27.200 ;
        RECT 7.000 27.100 7.300 28.200 ;
        RECT 9.400 27.500 9.800 29.900 ;
        RECT 10.200 27.700 10.600 29.900 ;
        RECT 12.300 29.200 12.900 29.900 ;
        RECT 12.300 28.900 13.000 29.200 ;
        RECT 14.600 28.900 15.000 29.900 ;
        RECT 16.800 29.200 17.200 29.900 ;
        RECT 16.800 28.900 17.800 29.200 ;
        RECT 12.600 28.500 13.000 28.900 ;
        RECT 14.700 28.600 15.000 28.900 ;
        RECT 14.700 28.300 16.100 28.600 ;
        RECT 15.700 28.200 16.100 28.300 ;
        RECT 16.600 28.200 17.000 28.600 ;
        RECT 17.400 28.500 17.800 28.900 ;
        RECT 11.700 27.700 12.100 27.800 ;
        RECT 10.200 27.400 12.100 27.700 ;
        RECT 8.600 27.100 9.400 27.200 ;
        RECT 3.900 26.800 9.400 27.100 ;
        RECT 3.000 26.400 3.400 26.500 ;
        RECT 1.500 26.100 3.400 26.400 ;
        RECT 1.500 26.000 1.900 26.100 ;
        RECT 2.300 25.700 2.700 25.800 ;
        RECT 0.600 25.400 2.700 25.700 ;
        RECT 0.600 21.100 1.000 25.400 ;
        RECT 3.900 25.200 4.200 26.800 ;
        RECT 7.500 26.700 7.900 26.800 ;
        RECT 7.000 26.200 7.400 26.300 ;
        RECT 8.300 26.200 8.700 26.300 ;
        RECT 6.200 25.900 8.700 26.200 ;
        RECT 6.200 25.800 6.600 25.900 ;
        RECT 10.200 25.700 10.600 27.400 ;
        RECT 13.700 27.100 14.100 27.200 ;
        RECT 16.600 27.100 16.900 28.200 ;
        RECT 19.000 27.500 19.400 29.900 ;
        RECT 19.800 27.500 20.200 29.900 ;
        RECT 22.000 29.200 22.400 29.900 ;
        RECT 21.400 28.900 22.400 29.200 ;
        RECT 24.200 28.900 24.600 29.900 ;
        RECT 26.300 29.200 26.900 29.900 ;
        RECT 26.200 28.900 26.900 29.200 ;
        RECT 21.400 28.500 21.800 28.900 ;
        RECT 24.200 28.600 24.500 28.900 ;
        RECT 22.200 28.200 22.600 28.600 ;
        RECT 23.100 28.300 24.500 28.600 ;
        RECT 26.200 28.500 26.600 28.900 ;
        RECT 23.100 28.200 23.500 28.300 ;
        RECT 18.200 27.100 19.000 27.200 ;
        RECT 20.200 27.100 21.000 27.200 ;
        RECT 22.300 27.100 22.600 28.200 ;
        RECT 27.100 27.700 27.500 27.800 ;
        RECT 28.600 27.700 29.000 29.900 ;
        RECT 30.700 28.200 31.100 29.900 ;
        RECT 27.100 27.400 29.000 27.700 ;
        RECT 30.200 27.900 31.100 28.200 ;
        RECT 25.100 27.100 25.800 27.200 ;
        RECT 13.500 26.800 25.800 27.100 ;
        RECT 28.600 27.100 29.000 27.400 ;
        RECT 29.400 27.100 29.800 27.600 ;
        RECT 28.600 26.800 29.800 27.100 ;
        RECT 12.600 26.400 13.000 26.500 ;
        RECT 11.100 26.100 13.000 26.400 ;
        RECT 13.500 26.200 13.800 26.800 ;
        RECT 17.100 26.700 17.500 26.800 ;
        RECT 21.700 26.700 22.100 26.800 ;
        RECT 16.600 26.200 17.000 26.300 ;
        RECT 17.900 26.200 18.300 26.300 ;
        RECT 11.100 26.000 11.500 26.100 ;
        RECT 13.400 25.800 13.800 26.200 ;
        RECT 15.800 25.900 18.300 26.200 ;
        RECT 20.900 26.200 21.300 26.300 ;
        RECT 20.900 25.900 23.400 26.200 ;
        RECT 15.800 25.800 16.200 25.900 ;
        RECT 23.000 25.800 23.400 25.900 ;
        RECT 11.900 25.700 12.300 25.800 ;
        RECT 7.000 25.500 9.800 25.600 ;
        RECT 6.900 25.400 9.800 25.500 ;
        RECT 3.000 24.900 4.200 25.200 ;
        RECT 4.900 25.300 9.800 25.400 ;
        RECT 4.900 25.100 7.300 25.300 ;
        RECT 3.000 24.400 3.300 24.900 ;
        RECT 2.600 24.000 3.300 24.400 ;
        RECT 4.100 24.500 4.500 24.600 ;
        RECT 4.900 24.500 5.200 25.100 ;
        RECT 4.100 24.200 5.200 24.500 ;
        RECT 5.500 24.500 8.200 24.800 ;
        RECT 5.500 24.400 5.900 24.500 ;
        RECT 7.800 24.400 8.200 24.500 ;
        RECT 4.700 23.700 5.100 23.800 ;
        RECT 6.100 23.700 6.500 23.800 ;
        RECT 3.000 23.100 3.400 23.500 ;
        RECT 4.700 23.400 6.500 23.700 ;
        RECT 5.100 23.100 5.400 23.400 ;
        RECT 7.800 23.100 8.200 23.500 ;
        RECT 2.700 21.100 3.300 23.100 ;
        RECT 5.000 21.100 5.400 23.100 ;
        RECT 7.200 22.800 8.200 23.100 ;
        RECT 7.200 21.100 7.600 22.800 ;
        RECT 9.400 21.100 9.800 25.300 ;
        RECT 10.200 25.400 12.300 25.700 ;
        RECT 10.200 21.100 10.600 25.400 ;
        RECT 13.500 25.200 13.800 25.800 ;
        RECT 16.600 25.500 19.400 25.600 ;
        RECT 16.500 25.400 19.400 25.500 ;
        RECT 12.600 24.900 13.800 25.200 ;
        RECT 14.500 25.300 19.400 25.400 ;
        RECT 14.500 25.100 16.900 25.300 ;
        RECT 12.600 24.400 12.900 24.900 ;
        RECT 12.200 24.000 12.900 24.400 ;
        RECT 13.700 24.500 14.100 24.600 ;
        RECT 14.500 24.500 14.800 25.100 ;
        RECT 13.700 24.200 14.800 24.500 ;
        RECT 15.100 24.500 17.800 24.800 ;
        RECT 15.100 24.400 15.500 24.500 ;
        RECT 17.400 24.400 17.800 24.500 ;
        RECT 14.300 23.700 14.700 23.800 ;
        RECT 15.700 23.700 16.100 23.800 ;
        RECT 12.600 23.100 13.000 23.500 ;
        RECT 14.300 23.400 16.100 23.700 ;
        RECT 14.700 23.100 15.000 23.400 ;
        RECT 17.400 23.100 17.800 23.500 ;
        RECT 12.300 21.100 12.900 23.100 ;
        RECT 14.600 21.100 15.000 23.100 ;
        RECT 16.800 22.800 17.800 23.100 ;
        RECT 16.800 21.100 17.200 22.800 ;
        RECT 19.000 21.100 19.400 25.300 ;
        RECT 19.800 25.500 22.600 25.600 ;
        RECT 19.800 25.400 22.700 25.500 ;
        RECT 19.800 25.300 24.700 25.400 ;
        RECT 19.800 21.100 20.200 25.300 ;
        RECT 22.300 25.100 24.700 25.300 ;
        RECT 21.400 24.500 24.100 24.800 ;
        RECT 21.400 24.400 21.800 24.500 ;
        RECT 23.700 24.400 24.100 24.500 ;
        RECT 24.400 24.500 24.700 25.100 ;
        RECT 25.400 25.200 25.700 26.800 ;
        RECT 26.200 26.400 26.600 26.500 ;
        RECT 26.200 26.100 28.100 26.400 ;
        RECT 27.700 26.000 28.100 26.100 ;
        RECT 26.900 25.700 27.300 25.800 ;
        RECT 28.600 25.700 29.000 26.800 ;
        RECT 26.900 25.400 29.000 25.700 ;
        RECT 25.400 24.900 26.600 25.200 ;
        RECT 25.100 24.500 25.500 24.600 ;
        RECT 24.400 24.200 25.500 24.500 ;
        RECT 26.300 24.400 26.600 24.900 ;
        RECT 26.300 24.000 27.000 24.400 ;
        RECT 23.100 23.700 23.500 23.800 ;
        RECT 24.500 23.700 24.900 23.800 ;
        RECT 21.400 23.100 21.800 23.500 ;
        RECT 23.100 23.400 24.900 23.700 ;
        RECT 24.200 23.100 24.500 23.400 ;
        RECT 26.200 23.100 26.600 23.500 ;
        RECT 21.400 22.800 22.400 23.100 ;
        RECT 22.000 21.100 22.400 22.800 ;
        RECT 24.200 21.100 24.600 23.100 ;
        RECT 26.300 21.100 26.900 23.100 ;
        RECT 28.600 21.100 29.000 25.400 ;
        RECT 30.200 26.100 30.600 27.900 ;
        RECT 31.800 27.800 32.200 29.900 ;
        RECT 32.600 28.000 33.000 29.900 ;
        RECT 34.200 28.000 34.600 29.900 ;
        RECT 32.600 27.900 34.600 28.000 ;
        RECT 31.900 27.200 32.200 27.800 ;
        RECT 32.700 27.700 34.500 27.900 ;
        RECT 35.000 27.500 35.400 29.900 ;
        RECT 37.200 29.200 37.600 29.900 ;
        RECT 36.600 28.900 37.600 29.200 ;
        RECT 39.400 28.900 39.800 29.900 ;
        RECT 41.500 29.200 42.100 29.900 ;
        RECT 41.400 28.900 42.100 29.200 ;
        RECT 36.600 28.500 37.000 28.900 ;
        RECT 39.400 28.600 39.700 28.900 ;
        RECT 37.400 28.200 37.800 28.600 ;
        RECT 38.300 28.300 39.700 28.600 ;
        RECT 41.400 28.500 41.800 28.900 ;
        RECT 38.300 28.200 38.700 28.300 ;
        RECT 33.800 27.200 34.200 27.400 ;
        RECT 31.800 26.800 33.100 27.200 ;
        RECT 33.800 26.900 34.600 27.200 ;
        RECT 34.200 26.800 34.600 26.900 ;
        RECT 35.400 27.100 36.200 27.200 ;
        RECT 37.500 27.100 37.800 28.200 ;
        RECT 42.300 27.700 42.700 27.800 ;
        RECT 43.800 27.700 44.200 29.900 ;
        RECT 44.600 28.000 45.000 29.900 ;
        RECT 46.200 28.000 46.600 29.900 ;
        RECT 44.600 27.900 46.600 28.000 ;
        RECT 47.000 27.900 47.400 29.900 ;
        RECT 48.100 28.200 48.500 29.900 ;
        RECT 52.600 28.200 53.000 29.900 ;
        RECT 48.100 27.900 49.000 28.200 ;
        RECT 44.700 27.700 46.500 27.900 ;
        RECT 42.300 27.400 44.200 27.700 ;
        RECT 40.300 27.100 40.700 27.200 ;
        RECT 35.400 26.800 40.900 27.100 ;
        RECT 30.200 25.800 32.100 26.100 ;
        RECT 30.200 21.100 30.600 25.800 ;
        RECT 31.800 25.200 32.100 25.800 ;
        RECT 31.000 24.400 31.400 25.200 ;
        RECT 31.800 25.100 32.200 25.200 ;
        RECT 32.800 25.100 33.100 26.800 ;
        RECT 36.900 26.700 37.300 26.800 ;
        RECT 33.400 25.800 33.800 26.600 ;
        RECT 36.100 26.200 36.500 26.300 ;
        RECT 36.100 25.900 38.600 26.200 ;
        RECT 38.200 25.800 38.600 25.900 ;
        RECT 35.000 25.500 37.800 25.600 ;
        RECT 35.000 25.400 37.900 25.500 ;
        RECT 35.000 25.300 39.900 25.400 ;
        RECT 31.800 24.800 32.500 25.100 ;
        RECT 32.800 24.800 33.300 25.100 ;
        RECT 32.200 24.200 32.500 24.800 ;
        RECT 32.200 23.800 32.600 24.200 ;
        RECT 32.900 21.100 33.300 24.800 ;
        RECT 35.000 21.100 35.400 25.300 ;
        RECT 37.500 25.100 39.900 25.300 ;
        RECT 36.600 24.500 39.300 24.800 ;
        RECT 36.600 24.400 37.000 24.500 ;
        RECT 38.900 24.400 39.300 24.500 ;
        RECT 39.600 24.500 39.900 25.100 ;
        RECT 40.600 25.200 40.900 26.800 ;
        RECT 41.400 26.400 41.800 26.500 ;
        RECT 41.400 26.100 43.300 26.400 ;
        RECT 42.900 26.000 43.300 26.100 ;
        RECT 42.100 25.700 42.500 25.800 ;
        RECT 43.800 25.700 44.200 27.400 ;
        RECT 45.000 27.200 45.400 27.400 ;
        RECT 47.000 27.200 47.300 27.900 ;
        RECT 44.600 26.900 45.400 27.200 ;
        RECT 44.600 26.800 45.000 26.900 ;
        RECT 46.100 26.800 47.400 27.200 ;
        RECT 45.400 25.800 45.800 26.600 ;
        RECT 42.100 25.400 44.200 25.700 ;
        RECT 40.600 24.900 41.800 25.200 ;
        RECT 40.300 24.500 40.700 24.600 ;
        RECT 39.600 24.200 40.700 24.500 ;
        RECT 41.500 24.400 41.800 24.900 ;
        RECT 41.500 24.000 42.200 24.400 ;
        RECT 38.300 23.700 38.700 23.800 ;
        RECT 39.700 23.700 40.100 23.800 ;
        RECT 36.600 23.100 37.000 23.500 ;
        RECT 38.300 23.400 40.100 23.700 ;
        RECT 39.400 23.100 39.700 23.400 ;
        RECT 41.400 23.100 41.800 23.500 ;
        RECT 36.600 22.800 37.600 23.100 ;
        RECT 37.200 21.100 37.600 22.800 ;
        RECT 39.400 21.100 39.800 23.100 ;
        RECT 41.500 21.100 42.100 23.100 ;
        RECT 43.800 21.100 44.200 25.400 ;
        RECT 46.100 25.200 46.400 26.800 ;
        RECT 48.600 26.100 49.000 27.900 ;
        RECT 52.500 27.900 53.000 28.200 ;
        RECT 49.400 26.800 49.800 27.600 ;
        RECT 52.500 27.200 52.800 27.900 ;
        RECT 54.200 27.600 54.600 29.900 ;
        RECT 55.000 28.000 55.400 29.900 ;
        RECT 56.600 28.000 57.000 29.900 ;
        RECT 55.000 27.900 57.000 28.000 ;
        RECT 57.400 28.100 57.800 29.900 ;
        RECT 58.300 28.200 58.700 28.600 ;
        RECT 58.200 28.100 58.600 28.200 ;
        RECT 55.100 27.700 56.900 27.900 ;
        RECT 57.400 27.800 58.600 28.100 ;
        RECT 59.000 27.900 59.400 29.900 ;
        RECT 62.200 28.900 62.600 29.900 ;
        RECT 53.300 27.300 54.600 27.600 ;
        RECT 50.200 27.100 50.600 27.200 ;
        RECT 52.500 27.100 53.000 27.200 ;
        RECT 50.200 26.800 53.000 27.100 ;
        RECT 45.400 24.800 46.400 25.200 ;
        RECT 47.000 25.800 49.000 26.100 ;
        RECT 47.000 25.200 47.300 25.800 ;
        RECT 47.000 25.100 47.400 25.200 ;
        RECT 46.700 24.800 47.400 25.100 ;
        RECT 45.900 21.100 46.300 24.800 ;
        RECT 46.700 24.200 47.000 24.800 ;
        RECT 47.800 24.400 48.200 25.200 ;
        RECT 46.600 23.800 47.000 24.200 ;
        RECT 48.600 21.100 49.000 25.800 ;
        RECT 52.500 25.100 52.800 26.800 ;
        RECT 53.300 26.500 53.600 27.300 ;
        RECT 55.400 27.200 55.800 27.400 ;
        RECT 57.400 27.200 57.700 27.800 ;
        RECT 55.000 26.900 55.800 27.200 ;
        RECT 55.000 26.800 55.400 26.900 ;
        RECT 56.500 26.800 57.800 27.200 ;
        RECT 53.100 26.100 53.600 26.500 ;
        RECT 53.300 25.100 53.600 26.100 ;
        RECT 54.100 26.200 54.500 26.600 ;
        RECT 54.100 25.800 54.600 26.200 ;
        RECT 55.800 25.800 56.200 26.600 ;
        RECT 56.500 25.100 56.800 26.800 ;
        RECT 58.200 26.100 58.600 26.200 ;
        RECT 59.100 26.100 59.400 27.900 ;
        RECT 61.400 27.800 61.800 28.600 ;
        RECT 62.300 28.100 62.600 28.900 ;
        RECT 62.200 27.800 63.300 28.100 ;
        RECT 63.800 27.900 64.200 29.900 ;
        RECT 64.600 28.000 65.000 29.900 ;
        RECT 66.200 28.000 66.600 29.900 ;
        RECT 64.600 27.900 66.600 28.000 ;
        RECT 67.000 28.000 67.400 29.900 ;
        RECT 68.600 28.000 69.000 29.900 ;
        RECT 67.000 27.900 69.000 28.000 ;
        RECT 69.400 27.900 69.800 29.900 ;
        RECT 70.200 27.900 70.600 29.900 ;
        RECT 71.000 28.000 71.400 29.900 ;
        RECT 72.600 28.000 73.000 29.900 ;
        RECT 75.300 29.200 75.700 29.500 ;
        RECT 75.000 28.800 75.700 29.200 ;
        RECT 75.300 28.000 75.700 28.800 ;
        RECT 77.400 28.500 77.800 29.500 ;
        RECT 71.000 27.900 73.000 28.000 ;
        RECT 62.300 27.200 62.600 27.800 ;
        RECT 59.800 26.400 60.200 27.200 ;
        RECT 62.200 26.800 62.600 27.200 ;
        RECT 63.000 27.200 63.300 27.800 ;
        RECT 63.900 27.200 64.200 27.900 ;
        RECT 64.700 27.700 66.500 27.900 ;
        RECT 67.100 27.700 68.900 27.900 ;
        RECT 65.800 27.200 66.200 27.400 ;
        RECT 67.400 27.200 67.800 27.400 ;
        RECT 69.400 27.200 69.700 27.900 ;
        RECT 70.300 27.200 70.600 27.900 ;
        RECT 71.100 27.700 72.900 27.900 ;
        RECT 74.900 27.700 75.700 28.000 ;
        RECT 74.900 27.500 75.300 27.700 ;
        RECT 72.200 27.200 72.600 27.400 ;
        RECT 74.900 27.200 75.200 27.500 ;
        RECT 77.500 27.400 77.800 28.500 ;
        RECT 79.500 28.200 79.900 29.900 ;
        RECT 79.000 27.900 79.900 28.200 ;
        RECT 80.600 27.900 81.000 29.900 ;
        RECT 81.400 28.000 81.800 29.900 ;
        RECT 83.000 28.000 83.400 29.900 ;
        RECT 81.400 27.900 83.400 28.000 ;
        RECT 83.800 28.000 84.200 29.900 ;
        RECT 85.400 28.000 85.800 29.900 ;
        RECT 83.800 27.900 85.800 28.000 ;
        RECT 86.200 27.900 86.600 29.900 ;
        RECT 87.000 28.500 87.400 29.500 ;
        RECT 63.000 26.800 63.400 27.200 ;
        RECT 63.800 26.800 65.100 27.200 ;
        RECT 65.800 26.900 66.600 27.200 ;
        RECT 66.200 26.800 66.600 26.900 ;
        RECT 67.000 26.900 67.800 27.200 ;
        RECT 67.000 26.800 67.400 26.900 ;
        RECT 68.500 26.800 69.800 27.200 ;
        RECT 70.200 26.800 71.500 27.200 ;
        RECT 72.200 26.900 73.000 27.200 ;
        RECT 72.600 26.800 73.000 26.900 ;
        RECT 74.200 26.800 75.200 27.200 ;
        RECT 75.700 27.100 77.800 27.400 ;
        RECT 75.700 26.900 76.200 27.100 ;
        RECT 60.600 26.100 61.000 26.200 ;
        RECT 58.200 25.800 59.400 26.100 ;
        RECT 60.200 25.800 61.000 26.100 ;
        RECT 57.400 25.100 57.800 25.200 ;
        RECT 58.300 25.100 58.600 25.800 ;
        RECT 60.200 25.600 60.600 25.800 ;
        RECT 62.300 25.100 62.600 26.800 ;
        RECT 63.000 25.400 63.400 26.200 ;
        RECT 64.800 25.200 65.100 26.800 ;
        RECT 65.400 26.100 65.800 26.600 ;
        RECT 66.200 26.100 66.600 26.200 ;
        RECT 65.400 25.800 66.600 26.100 ;
        RECT 67.800 25.800 68.200 26.600 ;
        RECT 63.800 25.100 64.200 25.200 ;
        RECT 52.500 24.600 53.000 25.100 ;
        RECT 53.300 24.800 54.600 25.100 ;
        RECT 52.600 21.100 53.000 24.600 ;
        RECT 54.200 21.100 54.600 24.800 ;
        RECT 56.300 24.800 56.800 25.100 ;
        RECT 57.100 24.800 57.800 25.100 ;
        RECT 56.300 21.100 56.700 24.800 ;
        RECT 57.100 24.200 57.400 24.800 ;
        RECT 57.000 23.800 57.400 24.200 ;
        RECT 58.200 21.100 58.600 25.100 ;
        RECT 59.000 24.800 61.000 25.100 ;
        RECT 59.000 21.100 59.400 24.800 ;
        RECT 60.600 21.100 61.000 24.800 ;
        RECT 62.200 24.700 63.100 25.100 ;
        RECT 63.800 24.800 64.500 25.100 ;
        RECT 64.800 24.800 65.800 25.200 ;
        RECT 68.500 25.100 68.800 26.800 ;
        RECT 71.200 25.200 71.500 26.800 ;
        RECT 71.800 26.100 72.200 26.600 ;
        RECT 72.600 26.100 73.000 26.200 ;
        RECT 71.800 25.800 73.000 26.100 ;
        RECT 74.200 25.400 74.600 26.200 ;
        RECT 69.400 25.100 69.800 25.200 ;
        RECT 68.300 24.800 68.800 25.100 ;
        RECT 69.100 24.800 69.800 25.100 ;
        RECT 70.200 25.100 70.600 25.200 ;
        RECT 70.200 24.800 70.900 25.100 ;
        RECT 71.200 24.800 72.200 25.200 ;
        RECT 74.900 24.900 75.200 26.800 ;
        RECT 75.500 26.500 76.200 26.900 ;
        RECT 78.200 26.800 78.600 27.600 ;
        RECT 75.900 25.500 76.200 26.500 ;
        RECT 76.600 25.800 77.000 26.600 ;
        RECT 77.400 25.800 77.800 26.600 ;
        RECT 79.000 26.100 79.400 27.900 ;
        RECT 80.700 27.200 81.000 27.900 ;
        RECT 81.500 27.700 83.300 27.900 ;
        RECT 83.900 27.700 85.700 27.900 ;
        RECT 82.600 27.200 83.000 27.400 ;
        RECT 84.200 27.200 84.600 27.400 ;
        RECT 86.200 27.200 86.500 27.900 ;
        RECT 87.000 27.400 87.300 28.500 ;
        RECT 89.100 28.000 89.500 29.500 ;
        RECT 91.800 28.000 92.200 29.900 ;
        RECT 93.400 28.000 93.800 29.900 ;
        RECT 89.100 27.700 89.900 28.000 ;
        RECT 91.800 27.900 93.800 28.000 ;
        RECT 94.200 27.900 94.600 29.900 ;
        RECT 95.000 28.000 95.400 29.900 ;
        RECT 96.600 28.000 97.000 29.900 ;
        RECT 95.000 27.900 97.000 28.000 ;
        RECT 97.400 27.900 97.800 29.900 ;
        RECT 98.200 28.500 98.600 29.500 ;
        RECT 91.900 27.700 93.700 27.900 ;
        RECT 89.500 27.500 89.900 27.700 ;
        RECT 80.600 26.800 81.900 27.200 ;
        RECT 82.600 26.900 83.400 27.200 ;
        RECT 83.000 26.800 83.400 26.900 ;
        RECT 83.800 26.900 84.600 27.200 ;
        RECT 83.800 26.800 84.200 26.900 ;
        RECT 85.300 26.800 86.600 27.200 ;
        RECT 87.000 27.100 89.100 27.400 ;
        RECT 88.600 26.900 89.100 27.100 ;
        RECT 89.600 27.200 89.900 27.500 ;
        RECT 92.200 27.200 92.600 27.400 ;
        RECT 94.200 27.200 94.500 27.900 ;
        RECT 95.100 27.700 96.900 27.900 ;
        RECT 95.400 27.200 95.800 27.400 ;
        RECT 97.400 27.200 97.700 27.900 ;
        RECT 98.200 27.400 98.500 28.500 ;
        RECT 100.300 28.000 100.700 29.500 ;
        RECT 104.700 28.200 105.100 28.600 ;
        RECT 100.300 27.700 101.100 28.000 ;
        RECT 104.600 27.800 105.000 28.200 ;
        RECT 105.400 27.900 105.800 29.900 ;
        RECT 108.600 28.900 109.000 29.900 ;
        RECT 100.700 27.500 101.100 27.700 ;
        RECT 81.600 26.200 81.900 26.800 ;
        RECT 79.000 25.800 80.900 26.100 ;
        RECT 81.400 25.800 81.900 26.200 ;
        RECT 82.200 25.800 82.600 26.600 ;
        RECT 83.000 26.100 83.400 26.200 ;
        RECT 84.600 26.100 85.000 26.600 ;
        RECT 83.000 25.800 85.000 26.100 ;
        RECT 75.900 25.200 77.800 25.500 ;
        RECT 62.700 21.100 63.100 24.700 ;
        RECT 64.200 24.200 64.500 24.800 ;
        RECT 64.200 23.800 64.600 24.200 ;
        RECT 64.900 21.100 65.300 24.800 ;
        RECT 68.300 21.100 68.700 24.800 ;
        RECT 69.100 24.200 69.400 24.800 ;
        RECT 69.000 23.800 69.400 24.200 ;
        RECT 70.600 24.200 70.900 24.800 ;
        RECT 70.600 23.800 71.000 24.200 ;
        RECT 71.300 21.100 71.700 24.800 ;
        RECT 74.900 24.600 75.700 24.900 ;
        RECT 75.300 21.100 75.700 24.600 ;
        RECT 77.500 23.500 77.800 25.200 ;
        RECT 77.400 21.500 77.800 23.500 ;
        RECT 79.000 21.100 79.400 25.800 ;
        RECT 80.600 25.200 80.900 25.800 ;
        RECT 79.800 24.400 80.200 25.200 ;
        RECT 80.600 25.100 81.000 25.200 ;
        RECT 81.600 25.100 81.900 25.800 ;
        RECT 85.300 25.100 85.600 26.800 ;
        RECT 87.000 25.800 87.400 26.600 ;
        RECT 87.800 25.800 88.200 26.600 ;
        RECT 88.600 26.500 89.300 26.900 ;
        RECT 89.600 26.800 90.600 27.200 ;
        RECT 91.800 26.900 92.600 27.200 ;
        RECT 91.800 26.800 92.200 26.900 ;
        RECT 93.300 26.800 94.600 27.200 ;
        RECT 95.000 26.900 95.800 27.200 ;
        RECT 95.000 26.800 95.400 26.900 ;
        RECT 96.500 26.800 97.800 27.200 ;
        RECT 98.200 27.100 100.300 27.400 ;
        RECT 99.800 26.900 100.300 27.100 ;
        RECT 100.800 27.200 101.100 27.500 ;
        RECT 88.600 25.500 88.900 26.500 ;
        RECT 87.000 25.200 88.900 25.500 ;
        RECT 86.200 25.100 86.600 25.200 ;
        RECT 80.600 24.800 81.300 25.100 ;
        RECT 81.600 24.800 82.100 25.100 ;
        RECT 81.000 24.200 81.300 24.800 ;
        RECT 81.000 23.800 81.400 24.200 ;
        RECT 81.700 21.100 82.100 24.800 ;
        RECT 85.100 24.800 85.600 25.100 ;
        RECT 85.900 24.800 86.600 25.100 ;
        RECT 85.100 21.100 85.500 24.800 ;
        RECT 85.900 24.200 86.200 24.800 ;
        RECT 85.800 23.800 86.200 24.200 ;
        RECT 87.000 23.500 87.300 25.200 ;
        RECT 89.600 24.900 89.900 26.800 ;
        RECT 90.200 25.400 90.600 26.200 ;
        RECT 92.600 25.800 93.000 26.600 ;
        RECT 93.300 25.100 93.600 26.800 ;
        RECT 95.800 25.800 96.200 26.600 ;
        RECT 96.500 26.100 96.800 26.800 ;
        RECT 97.400 26.100 97.800 26.200 ;
        RECT 96.500 25.800 97.800 26.100 ;
        RECT 98.200 25.800 98.600 26.600 ;
        RECT 99.000 25.800 99.400 26.600 ;
        RECT 99.800 26.500 100.500 26.900 ;
        RECT 100.800 26.800 101.800 27.200 ;
        RECT 94.200 25.100 94.600 25.200 ;
        RECT 96.500 25.100 96.800 25.800 ;
        RECT 99.800 25.500 100.100 26.500 ;
        RECT 98.200 25.200 100.100 25.500 ;
        RECT 97.400 25.100 97.800 25.200 ;
        RECT 89.100 24.600 89.900 24.900 ;
        RECT 93.100 24.800 93.600 25.100 ;
        RECT 93.900 24.800 94.600 25.100 ;
        RECT 96.300 24.800 96.800 25.100 ;
        RECT 97.100 24.800 97.800 25.100 ;
        RECT 87.000 21.500 87.400 23.500 ;
        RECT 89.100 22.200 89.500 24.600 ;
        RECT 89.100 21.800 89.800 22.200 ;
        RECT 89.100 21.100 89.500 21.800 ;
        RECT 93.100 21.100 93.500 24.800 ;
        RECT 93.900 24.200 94.200 24.800 ;
        RECT 93.800 23.800 94.200 24.200 ;
        RECT 96.300 21.100 96.700 24.800 ;
        RECT 97.100 24.200 97.400 24.800 ;
        RECT 97.000 23.800 97.400 24.200 ;
        RECT 98.200 23.500 98.500 25.200 ;
        RECT 100.800 24.900 101.100 26.800 ;
        RECT 101.400 25.400 101.800 26.200 ;
        RECT 104.600 26.100 105.000 26.200 ;
        RECT 105.500 26.100 105.800 27.900 ;
        RECT 107.800 27.800 108.200 28.600 ;
        RECT 108.700 28.100 109.000 28.900 ;
        RECT 110.300 28.200 110.700 28.600 ;
        RECT 110.200 28.100 110.600 28.200 ;
        RECT 108.600 27.800 110.600 28.100 ;
        RECT 111.000 27.900 111.400 29.900 ;
        RECT 113.400 27.900 113.800 29.900 ;
        RECT 114.200 28.000 114.600 29.900 ;
        RECT 115.800 28.000 116.200 29.900 ;
        RECT 114.200 27.900 116.200 28.000 ;
        RECT 116.600 27.900 117.000 29.900 ;
        RECT 117.400 28.000 117.800 29.900 ;
        RECT 119.000 28.000 119.400 29.900 ;
        RECT 117.400 27.900 119.400 28.000 ;
        RECT 119.800 27.900 120.200 29.900 ;
        RECT 120.600 28.000 121.000 29.900 ;
        RECT 122.200 28.000 122.600 29.900 ;
        RECT 120.600 27.900 122.600 28.000 ;
        RECT 123.000 28.000 123.400 29.900 ;
        RECT 124.600 28.000 125.000 29.900 ;
        RECT 123.000 27.900 125.000 28.000 ;
        RECT 125.400 27.900 125.800 29.900 ;
        RECT 127.800 27.900 128.200 29.900 ;
        RECT 128.500 28.200 128.900 28.600 ;
        RECT 128.600 28.100 129.000 28.200 ;
        RECT 129.400 28.100 129.800 29.900 ;
        RECT 106.200 27.100 106.600 27.200 ;
        RECT 107.800 27.100 108.100 27.800 ;
        RECT 108.700 27.200 109.000 27.800 ;
        RECT 106.200 26.800 108.100 27.100 ;
        RECT 108.600 26.800 109.000 27.200 ;
        RECT 106.200 26.400 106.600 26.800 ;
        RECT 107.000 26.100 107.400 26.200 ;
        RECT 104.600 25.800 105.800 26.100 ;
        RECT 106.600 25.800 107.400 26.100 ;
        RECT 104.700 25.100 105.000 25.800 ;
        RECT 106.600 25.600 107.000 25.800 ;
        RECT 108.700 25.100 109.000 26.800 ;
        RECT 109.400 25.400 109.800 26.200 ;
        RECT 110.200 26.100 110.600 26.200 ;
        RECT 111.100 26.100 111.400 27.900 ;
        RECT 113.500 27.200 113.800 27.900 ;
        RECT 114.300 27.700 116.100 27.900 ;
        RECT 115.400 27.200 115.800 27.400 ;
        RECT 116.700 27.200 117.000 27.900 ;
        RECT 117.500 27.700 119.300 27.900 ;
        RECT 118.600 27.200 119.000 27.400 ;
        RECT 119.900 27.200 120.200 27.900 ;
        RECT 120.700 27.700 122.500 27.900 ;
        RECT 123.100 27.700 124.900 27.900 ;
        RECT 121.800 27.200 122.200 27.400 ;
        RECT 123.400 27.200 123.800 27.400 ;
        RECT 125.400 27.200 125.700 27.900 ;
        RECT 111.800 26.400 112.200 27.200 ;
        RECT 112.600 27.100 113.000 27.200 ;
        RECT 113.400 27.100 114.700 27.200 ;
        RECT 112.600 26.800 114.700 27.100 ;
        RECT 115.400 26.900 116.200 27.200 ;
        RECT 115.800 26.800 116.200 26.900 ;
        RECT 116.600 26.800 117.900 27.200 ;
        RECT 118.600 26.900 119.400 27.200 ;
        RECT 119.000 26.800 119.400 26.900 ;
        RECT 119.800 26.800 121.100 27.200 ;
        RECT 121.800 27.100 122.600 27.200 ;
        RECT 123.000 27.100 123.800 27.200 ;
        RECT 121.800 26.900 123.800 27.100 ;
        RECT 122.200 26.800 123.400 26.900 ;
        RECT 124.500 26.800 125.800 27.200 ;
        RECT 112.600 26.100 113.000 26.200 ;
        RECT 110.200 25.800 111.400 26.100 ;
        RECT 112.200 25.800 113.000 26.100 ;
        RECT 110.300 25.100 110.600 25.800 ;
        RECT 112.200 25.600 112.600 25.800 ;
        RECT 113.400 25.100 113.800 25.200 ;
        RECT 114.400 25.100 114.700 26.800 ;
        RECT 115.000 25.800 115.400 26.600 ;
        RECT 116.600 25.100 117.000 25.200 ;
        RECT 117.600 25.100 117.900 26.800 ;
        RECT 118.200 26.100 118.600 26.600 ;
        RECT 119.000 26.100 119.400 26.200 ;
        RECT 118.200 25.800 119.400 26.100 ;
        RECT 119.800 26.100 120.200 26.200 ;
        RECT 120.800 26.100 121.100 26.800 ;
        RECT 119.800 25.800 121.100 26.100 ;
        RECT 121.400 25.800 121.800 26.600 ;
        RECT 123.800 25.800 124.200 26.600 ;
        RECT 119.800 25.100 120.200 25.200 ;
        RECT 120.800 25.100 121.100 25.800 ;
        RECT 124.500 25.100 124.800 26.800 ;
        RECT 127.000 26.400 127.400 27.200 ;
        RECT 126.200 26.100 126.600 26.200 ;
        RECT 127.800 26.100 128.100 27.900 ;
        RECT 128.600 27.800 129.800 28.100 ;
        RECT 130.200 28.000 130.600 29.900 ;
        RECT 131.800 28.000 132.200 29.900 ;
        RECT 130.200 27.900 132.200 28.000 ;
        RECT 129.500 27.200 129.800 27.800 ;
        RECT 130.300 27.700 132.100 27.900 ;
        RECT 132.600 27.700 133.000 29.900 ;
        RECT 134.700 29.200 135.300 29.900 ;
        RECT 134.700 28.900 135.400 29.200 ;
        RECT 137.000 28.900 137.400 29.900 ;
        RECT 139.200 29.200 139.600 29.900 ;
        RECT 139.200 28.900 140.200 29.200 ;
        RECT 135.000 28.500 135.400 28.900 ;
        RECT 137.100 28.600 137.400 28.900 ;
        RECT 137.100 28.300 138.500 28.600 ;
        RECT 138.100 28.200 138.500 28.300 ;
        RECT 139.000 28.200 139.400 28.600 ;
        RECT 139.800 28.500 140.200 28.900 ;
        RECT 134.100 27.700 134.500 27.800 ;
        RECT 132.600 27.400 134.500 27.700 ;
        RECT 131.400 27.200 131.800 27.400 ;
        RECT 129.400 26.800 130.700 27.200 ;
        RECT 131.400 26.900 132.200 27.200 ;
        RECT 131.800 26.800 132.200 26.900 ;
        RECT 128.600 26.100 129.000 26.200 ;
        RECT 126.200 25.800 127.000 26.100 ;
        RECT 127.800 25.800 129.000 26.100 ;
        RECT 126.600 25.600 127.000 25.800 ;
        RECT 125.400 25.100 125.800 25.200 ;
        RECT 128.600 25.100 128.900 25.800 ;
        RECT 129.400 25.100 129.800 25.200 ;
        RECT 130.400 25.100 130.700 26.800 ;
        RECT 131.000 25.800 131.400 26.600 ;
        RECT 132.600 25.700 133.000 27.400 ;
        RECT 136.100 27.100 136.500 27.200 ;
        RECT 139.000 27.100 139.300 28.200 ;
        RECT 141.400 27.500 141.800 29.900 ;
        RECT 143.000 28.800 143.400 29.900 ;
        RECT 142.200 27.800 142.600 28.600 ;
        RECT 143.100 27.200 143.400 28.800 ;
        RECT 140.600 27.100 141.400 27.200 ;
        RECT 135.900 26.800 141.400 27.100 ;
        RECT 143.000 26.800 143.400 27.200 ;
        RECT 135.000 26.400 135.400 26.500 ;
        RECT 133.500 26.100 135.400 26.400 ;
        RECT 133.500 26.000 133.900 26.100 ;
        RECT 134.300 25.700 134.700 25.800 ;
        RECT 132.600 25.400 134.700 25.700 ;
        RECT 100.300 24.600 101.100 24.900 ;
        RECT 98.200 21.500 98.600 23.500 ;
        RECT 100.300 22.200 100.700 24.600 ;
        RECT 100.300 21.800 101.000 22.200 ;
        RECT 100.300 21.100 100.700 21.800 ;
        RECT 104.600 21.100 105.000 25.100 ;
        RECT 105.400 24.800 107.400 25.100 ;
        RECT 105.400 21.100 105.800 24.800 ;
        RECT 107.000 21.100 107.400 24.800 ;
        RECT 108.600 24.700 109.500 25.100 ;
        RECT 109.100 21.100 109.500 24.700 ;
        RECT 110.200 21.100 110.600 25.100 ;
        RECT 111.000 24.800 113.000 25.100 ;
        RECT 113.400 24.800 114.100 25.100 ;
        RECT 114.400 24.800 114.900 25.100 ;
        RECT 116.600 24.800 117.300 25.100 ;
        RECT 117.600 24.800 118.100 25.100 ;
        RECT 119.800 24.800 120.500 25.100 ;
        RECT 120.800 24.800 121.300 25.100 ;
        RECT 111.000 21.100 111.400 24.800 ;
        RECT 112.600 21.100 113.000 24.800 ;
        RECT 113.800 24.200 114.100 24.800 ;
        RECT 113.800 23.800 114.200 24.200 ;
        RECT 114.500 21.100 114.900 24.800 ;
        RECT 117.000 24.200 117.300 24.800 ;
        RECT 117.000 23.800 117.400 24.200 ;
        RECT 117.700 22.200 118.100 24.800 ;
        RECT 120.200 24.200 120.500 24.800 ;
        RECT 120.200 23.800 120.600 24.200 ;
        RECT 117.700 21.800 118.600 22.200 ;
        RECT 117.700 21.100 118.100 21.800 ;
        RECT 120.900 21.100 121.300 24.800 ;
        RECT 124.300 24.800 124.800 25.100 ;
        RECT 125.100 24.800 125.800 25.100 ;
        RECT 126.200 24.800 128.200 25.100 ;
        RECT 124.300 21.100 124.700 24.800 ;
        RECT 125.100 24.200 125.400 24.800 ;
        RECT 125.000 23.800 125.400 24.200 ;
        RECT 126.200 21.100 126.600 24.800 ;
        RECT 127.800 21.100 128.200 24.800 ;
        RECT 128.600 21.100 129.000 25.100 ;
        RECT 129.400 24.800 130.100 25.100 ;
        RECT 130.400 24.800 130.900 25.100 ;
        RECT 129.800 24.200 130.100 24.800 ;
        RECT 129.800 23.800 130.200 24.200 ;
        RECT 130.500 21.100 130.900 24.800 ;
        RECT 132.600 21.100 133.000 25.400 ;
        RECT 135.900 25.200 136.200 26.800 ;
        RECT 139.500 26.700 139.900 26.800 ;
        RECT 140.300 26.200 140.700 26.300 ;
        RECT 136.600 26.100 137.000 26.200 ;
        RECT 138.200 26.100 140.700 26.200 ;
        RECT 136.600 25.900 140.700 26.100 ;
        RECT 136.600 25.800 138.600 25.900 ;
        RECT 139.000 25.500 141.800 25.600 ;
        RECT 138.900 25.400 141.800 25.500 ;
        RECT 135.000 24.900 136.200 25.200 ;
        RECT 136.900 25.300 141.800 25.400 ;
        RECT 136.900 25.100 139.300 25.300 ;
        RECT 135.000 24.400 135.300 24.900 ;
        RECT 134.600 24.000 135.300 24.400 ;
        RECT 136.100 24.500 136.500 24.600 ;
        RECT 136.900 24.500 137.200 25.100 ;
        RECT 136.100 24.200 137.200 24.500 ;
        RECT 137.500 24.500 140.200 24.800 ;
        RECT 137.500 24.400 137.900 24.500 ;
        RECT 139.800 24.400 140.200 24.500 ;
        RECT 136.700 23.700 137.100 23.800 ;
        RECT 138.100 23.700 138.500 23.800 ;
        RECT 135.000 23.100 135.400 23.500 ;
        RECT 136.700 23.400 138.500 23.700 ;
        RECT 137.100 23.100 137.400 23.400 ;
        RECT 139.800 23.100 140.200 23.500 ;
        RECT 134.700 21.100 135.300 23.100 ;
        RECT 137.000 21.100 137.400 23.100 ;
        RECT 139.200 22.800 140.200 23.100 ;
        RECT 139.200 21.100 139.600 22.800 ;
        RECT 141.400 21.100 141.800 25.300 ;
        RECT 143.100 25.100 143.400 26.800 ;
        RECT 144.600 27.700 145.000 29.900 ;
        RECT 146.700 29.200 147.300 29.900 ;
        RECT 146.700 28.900 147.400 29.200 ;
        RECT 149.000 28.900 149.400 29.900 ;
        RECT 151.200 29.200 151.600 29.900 ;
        RECT 151.200 28.900 152.200 29.200 ;
        RECT 147.000 28.500 147.400 28.900 ;
        RECT 149.100 28.600 149.400 28.900 ;
        RECT 149.100 28.300 150.500 28.600 ;
        RECT 150.100 28.200 150.500 28.300 ;
        RECT 151.000 28.200 151.400 28.600 ;
        RECT 151.800 28.500 152.200 28.900 ;
        RECT 146.100 27.700 146.500 27.800 ;
        RECT 144.600 27.400 146.500 27.700 ;
        RECT 143.800 25.400 144.200 26.200 ;
        RECT 144.600 25.700 145.000 27.400 ;
        RECT 148.100 27.100 148.500 27.200 ;
        RECT 151.000 27.100 151.300 28.200 ;
        RECT 153.400 27.500 153.800 29.900 ;
        RECT 157.400 27.900 157.800 29.900 ;
        RECT 159.800 28.900 160.200 29.900 ;
        RECT 158.100 28.200 158.500 28.600 ;
        RECT 152.600 27.100 153.400 27.200 ;
        RECT 147.900 26.800 153.400 27.100 ;
        RECT 147.000 26.400 147.400 26.500 ;
        RECT 145.500 26.100 147.400 26.400 ;
        RECT 147.900 26.100 148.200 26.800 ;
        RECT 151.500 26.700 151.900 26.800 ;
        RECT 156.600 26.400 157.000 27.200 ;
        RECT 151.000 26.200 151.400 26.300 ;
        RECT 152.300 26.200 152.700 26.300 ;
        RECT 148.600 26.100 149.000 26.200 ;
        RECT 145.500 26.000 145.900 26.100 ;
        RECT 147.800 25.800 149.000 26.100 ;
        RECT 150.200 25.900 152.700 26.200 ;
        RECT 154.200 26.100 154.600 26.200 ;
        RECT 155.800 26.100 156.200 26.200 ;
        RECT 157.400 26.100 157.700 27.900 ;
        RECT 158.200 27.800 158.600 28.200 ;
        RECT 159.000 27.800 159.400 28.600 ;
        RECT 158.200 27.100 158.500 27.800 ;
        RECT 159.900 27.200 160.200 28.900 ;
        RECT 161.500 28.200 161.900 28.600 ;
        RECT 161.400 27.800 161.800 28.200 ;
        RECT 162.200 27.900 162.600 29.900 ;
        RECT 164.600 27.900 165.000 29.900 ;
        RECT 165.400 28.000 165.800 29.900 ;
        RECT 167.000 28.000 167.400 29.900 ;
        RECT 165.400 27.900 167.400 28.000 ;
        RECT 159.800 27.100 160.200 27.200 ;
        RECT 158.200 26.800 160.200 27.100 ;
        RECT 158.200 26.100 158.600 26.200 ;
        RECT 150.200 25.800 150.600 25.900 ;
        RECT 154.200 25.800 156.600 26.100 ;
        RECT 157.400 25.800 158.600 26.100 ;
        RECT 146.300 25.700 146.700 25.800 ;
        RECT 144.600 25.400 146.700 25.700 ;
        RECT 143.000 24.700 143.900 25.100 ;
        RECT 143.500 21.100 143.900 24.700 ;
        RECT 144.600 21.100 145.000 25.400 ;
        RECT 147.900 25.200 148.200 25.800 ;
        RECT 156.200 25.600 156.600 25.800 ;
        RECT 151.000 25.500 153.800 25.600 ;
        RECT 150.900 25.400 153.800 25.500 ;
        RECT 147.000 24.900 148.200 25.200 ;
        RECT 148.900 25.300 153.800 25.400 ;
        RECT 148.900 25.100 151.300 25.300 ;
        RECT 147.000 24.400 147.300 24.900 ;
        RECT 146.600 24.200 147.300 24.400 ;
        RECT 148.100 24.500 148.500 24.600 ;
        RECT 148.900 24.500 149.200 25.100 ;
        RECT 148.100 24.200 149.200 24.500 ;
        RECT 149.500 24.500 152.200 24.800 ;
        RECT 149.500 24.400 149.900 24.500 ;
        RECT 151.800 24.400 152.200 24.500 ;
        RECT 146.200 24.000 147.300 24.200 ;
        RECT 146.200 23.800 146.900 24.000 ;
        RECT 148.700 23.700 149.100 23.800 ;
        RECT 150.100 23.700 150.500 23.800 ;
        RECT 147.000 23.100 147.400 23.500 ;
        RECT 148.700 23.400 150.500 23.700 ;
        RECT 149.100 23.100 149.400 23.400 ;
        RECT 151.800 23.100 152.200 23.500 ;
        RECT 146.700 21.100 147.300 23.100 ;
        RECT 149.000 21.100 149.400 23.100 ;
        RECT 151.200 22.800 152.200 23.100 ;
        RECT 151.200 21.100 151.600 22.800 ;
        RECT 153.400 21.100 153.800 25.300 ;
        RECT 158.200 25.100 158.500 25.800 ;
        RECT 159.900 25.100 160.200 26.800 ;
        RECT 162.300 26.200 162.600 27.900 ;
        RECT 164.700 27.200 165.000 27.900 ;
        RECT 165.500 27.700 167.300 27.900 ;
        RECT 167.800 27.700 168.200 29.900 ;
        RECT 169.900 29.200 170.500 29.900 ;
        RECT 169.900 28.900 170.600 29.200 ;
        RECT 172.200 28.900 172.600 29.900 ;
        RECT 174.400 29.200 174.800 29.900 ;
        RECT 174.400 28.900 175.400 29.200 ;
        RECT 170.200 28.500 170.600 28.900 ;
        RECT 172.300 28.600 172.600 28.900 ;
        RECT 172.300 28.300 173.700 28.600 ;
        RECT 173.300 28.200 173.700 28.300 ;
        RECT 174.200 28.200 174.600 28.600 ;
        RECT 175.000 28.500 175.400 28.900 ;
        RECT 169.300 27.700 169.700 27.800 ;
        RECT 167.800 27.400 169.700 27.700 ;
        RECT 166.600 27.200 167.000 27.400 ;
        RECT 163.000 26.400 163.400 27.200 ;
        RECT 164.600 26.800 165.900 27.200 ;
        RECT 166.600 26.900 167.400 27.200 ;
        RECT 167.000 26.800 167.400 26.900 ;
        RECT 160.600 25.400 161.000 26.200 ;
        RECT 161.400 26.100 161.800 26.200 ;
        RECT 162.200 26.100 162.600 26.200 ;
        RECT 163.800 26.100 164.200 26.200 ;
        RECT 161.400 25.800 162.600 26.100 ;
        RECT 163.400 25.800 164.200 26.100 ;
        RECT 161.500 25.100 161.800 25.800 ;
        RECT 163.400 25.600 163.800 25.800 ;
        RECT 164.600 25.100 165.000 25.200 ;
        RECT 165.600 25.100 165.900 26.800 ;
        RECT 166.200 26.100 166.600 26.600 ;
        RECT 167.000 26.100 167.400 26.200 ;
        RECT 166.200 25.800 167.400 26.100 ;
        RECT 167.800 25.700 168.200 27.400 ;
        RECT 171.300 27.100 171.700 27.200 ;
        RECT 174.200 27.100 174.500 28.200 ;
        RECT 176.600 27.500 177.000 29.900 ;
        RECT 177.400 27.700 177.800 29.900 ;
        RECT 179.500 29.200 180.100 29.900 ;
        RECT 179.500 28.900 180.200 29.200 ;
        RECT 181.800 28.900 182.200 29.900 ;
        RECT 184.000 29.200 184.400 29.900 ;
        RECT 184.000 28.900 185.000 29.200 ;
        RECT 179.800 28.500 180.200 28.900 ;
        RECT 181.900 28.600 182.200 28.900 ;
        RECT 181.900 28.300 183.300 28.600 ;
        RECT 182.900 28.200 183.300 28.300 ;
        RECT 183.800 28.200 184.200 28.600 ;
        RECT 184.600 28.500 185.000 28.900 ;
        RECT 179.000 27.800 179.400 28.200 ;
        RECT 178.900 27.700 179.400 27.800 ;
        RECT 177.400 27.400 179.400 27.700 ;
        RECT 175.800 27.100 176.600 27.200 ;
        RECT 171.100 26.800 176.600 27.100 ;
        RECT 170.200 26.400 170.600 26.500 ;
        RECT 168.700 26.100 170.600 26.400 ;
        RECT 168.700 26.000 169.100 26.100 ;
        RECT 169.500 25.700 169.900 25.800 ;
        RECT 167.800 25.400 169.900 25.700 ;
        RECT 155.800 24.800 157.800 25.100 ;
        RECT 155.800 21.100 156.200 24.800 ;
        RECT 157.400 21.100 157.800 24.800 ;
        RECT 158.200 21.100 158.600 25.100 ;
        RECT 159.800 24.700 160.700 25.100 ;
        RECT 160.300 21.100 160.700 24.700 ;
        RECT 161.400 21.100 161.800 25.100 ;
        RECT 162.200 24.800 164.200 25.100 ;
        RECT 164.600 24.800 165.300 25.100 ;
        RECT 165.600 24.800 166.100 25.100 ;
        RECT 162.200 21.100 162.600 24.800 ;
        RECT 163.800 21.100 164.200 24.800 ;
        RECT 165.000 24.200 165.300 24.800 ;
        RECT 165.000 23.800 165.400 24.200 ;
        RECT 165.700 21.100 166.100 24.800 ;
        RECT 167.800 21.100 168.200 25.400 ;
        RECT 171.100 25.200 171.400 26.800 ;
        RECT 174.700 26.700 175.100 26.800 ;
        RECT 175.500 26.200 175.900 26.300 ;
        RECT 171.800 26.100 172.200 26.200 ;
        RECT 173.400 26.100 175.900 26.200 ;
        RECT 171.800 25.900 175.900 26.100 ;
        RECT 171.800 25.800 173.800 25.900 ;
        RECT 177.400 25.700 177.800 27.400 ;
        RECT 180.900 27.100 181.300 27.200 ;
        RECT 183.800 27.100 184.100 28.200 ;
        RECT 186.200 27.500 186.600 29.900 ;
        RECT 187.000 28.500 187.400 29.500 ;
        RECT 187.000 27.400 187.300 28.500 ;
        RECT 189.100 28.000 189.500 29.500 ;
        RECT 189.100 27.700 189.900 28.000 ;
        RECT 189.500 27.500 189.900 27.700 ;
        RECT 185.400 27.100 186.200 27.200 ;
        RECT 187.000 27.100 189.100 27.400 ;
        RECT 180.700 26.800 186.200 27.100 ;
        RECT 188.600 26.900 189.100 27.100 ;
        RECT 189.600 27.200 189.900 27.500 ;
        RECT 179.800 26.400 180.200 26.500 ;
        RECT 178.300 26.100 180.200 26.400 ;
        RECT 180.700 26.200 181.000 26.800 ;
        RECT 184.300 26.700 184.700 26.800 ;
        RECT 185.100 26.200 185.500 26.300 ;
        RECT 178.300 26.000 178.700 26.100 ;
        RECT 180.600 25.800 181.000 26.200 ;
        RECT 183.000 25.900 185.500 26.200 ;
        RECT 183.000 25.800 183.400 25.900 ;
        RECT 187.000 25.800 187.400 26.600 ;
        RECT 187.800 25.800 188.200 26.600 ;
        RECT 188.600 26.500 189.300 26.900 ;
        RECT 189.600 26.800 190.600 27.200 ;
        RECT 179.100 25.700 179.500 25.800 ;
        RECT 174.200 25.500 177.000 25.600 ;
        RECT 174.100 25.400 177.000 25.500 ;
        RECT 170.200 24.900 171.400 25.200 ;
        RECT 172.100 25.300 177.000 25.400 ;
        RECT 172.100 25.100 174.500 25.300 ;
        RECT 170.200 24.400 170.500 24.900 ;
        RECT 169.800 24.200 170.500 24.400 ;
        RECT 171.300 24.500 171.700 24.600 ;
        RECT 172.100 24.500 172.400 25.100 ;
        RECT 171.300 24.200 172.400 24.500 ;
        RECT 172.700 24.500 175.400 24.800 ;
        RECT 172.700 24.400 173.100 24.500 ;
        RECT 175.000 24.400 175.400 24.500 ;
        RECT 169.400 24.000 170.500 24.200 ;
        RECT 169.400 23.800 170.100 24.000 ;
        RECT 171.900 23.700 172.300 23.800 ;
        RECT 173.300 23.700 173.700 23.800 ;
        RECT 170.200 23.100 170.600 23.500 ;
        RECT 171.900 23.400 173.700 23.700 ;
        RECT 172.300 23.100 172.600 23.400 ;
        RECT 175.000 23.100 175.400 23.500 ;
        RECT 169.900 21.100 170.500 23.100 ;
        RECT 172.200 21.100 172.600 23.100 ;
        RECT 174.400 22.800 175.400 23.100 ;
        RECT 174.400 21.100 174.800 22.800 ;
        RECT 176.600 21.100 177.000 25.300 ;
        RECT 177.400 25.400 179.500 25.700 ;
        RECT 177.400 21.100 177.800 25.400 ;
        RECT 180.700 25.200 181.000 25.800 ;
        RECT 183.800 25.500 186.600 25.600 ;
        RECT 188.600 25.500 188.900 26.500 ;
        RECT 183.700 25.400 186.600 25.500 ;
        RECT 179.800 24.900 181.000 25.200 ;
        RECT 181.700 25.300 186.600 25.400 ;
        RECT 181.700 25.100 184.100 25.300 ;
        RECT 179.800 24.400 180.100 24.900 ;
        RECT 179.400 24.000 180.100 24.400 ;
        RECT 180.900 24.500 181.300 24.600 ;
        RECT 181.700 24.500 182.000 25.100 ;
        RECT 180.900 24.200 182.000 24.500 ;
        RECT 182.300 24.500 185.000 24.800 ;
        RECT 182.300 24.400 182.700 24.500 ;
        RECT 184.600 24.400 185.000 24.500 ;
        RECT 181.500 23.700 181.900 23.800 ;
        RECT 182.900 23.700 183.300 23.800 ;
        RECT 179.800 23.100 180.200 23.500 ;
        RECT 181.500 23.400 183.300 23.700 ;
        RECT 181.900 23.100 182.200 23.400 ;
        RECT 184.600 23.100 185.000 23.500 ;
        RECT 179.500 21.100 180.100 23.100 ;
        RECT 181.800 21.100 182.200 23.100 ;
        RECT 184.000 22.800 185.000 23.100 ;
        RECT 184.000 21.100 184.400 22.800 ;
        RECT 186.200 21.100 186.600 25.300 ;
        RECT 187.000 25.200 188.900 25.500 ;
        RECT 187.000 23.500 187.300 25.200 ;
        RECT 189.600 24.900 189.900 26.800 ;
        RECT 190.200 25.400 190.600 26.200 ;
        RECT 189.100 24.600 189.900 24.900 ;
        RECT 187.000 21.500 187.400 23.500 ;
        RECT 189.100 22.200 189.500 24.600 ;
        RECT 189.100 21.800 189.800 22.200 ;
        RECT 189.100 21.100 189.500 21.800 ;
        RECT 191.800 21.100 192.200 29.900 ;
        RECT 192.600 26.800 193.000 27.600 ;
        RECT 193.400 21.100 193.800 29.900 ;
        RECT 194.200 27.800 194.600 28.600 ;
        RECT 195.000 28.500 195.400 29.500 ;
        RECT 195.000 27.400 195.300 28.500 ;
        RECT 197.100 28.000 197.500 29.500 ;
        RECT 197.100 27.700 197.900 28.000 ;
        RECT 197.500 27.500 197.900 27.700 ;
        RECT 201.400 27.600 201.800 29.900 ;
        RECT 195.000 27.100 197.100 27.400 ;
        RECT 196.600 26.900 197.100 27.100 ;
        RECT 197.600 27.200 197.900 27.500 ;
        RECT 200.700 27.300 201.800 27.600 ;
        RECT 202.200 27.600 202.600 29.900 ;
        RECT 202.200 27.300 203.300 27.600 ;
        RECT 194.200 26.100 194.600 26.200 ;
        RECT 195.000 26.100 195.400 26.600 ;
        RECT 194.200 25.800 195.400 26.100 ;
        RECT 195.800 25.800 196.200 26.600 ;
        RECT 196.600 26.500 197.300 26.900 ;
        RECT 197.600 26.800 198.600 27.200 ;
        RECT 196.600 25.500 196.900 26.500 ;
        RECT 195.000 25.200 196.900 25.500 ;
        RECT 195.000 23.500 195.300 25.200 ;
        RECT 197.600 24.900 197.900 26.800 ;
        RECT 198.200 25.400 198.600 26.200 ;
        RECT 200.700 25.800 201.000 27.300 ;
        RECT 201.400 25.800 201.800 26.600 ;
        RECT 202.200 25.800 202.600 26.600 ;
        RECT 203.000 25.800 203.300 27.300 ;
        RECT 200.400 25.400 201.000 25.800 ;
        RECT 197.100 24.600 197.900 24.900 ;
        RECT 200.700 25.100 201.000 25.400 ;
        RECT 203.000 25.400 203.600 25.800 ;
        RECT 203.000 25.100 203.300 25.400 ;
        RECT 200.700 24.800 201.800 25.100 ;
        RECT 195.000 21.500 195.400 23.500 ;
        RECT 197.100 22.200 197.500 24.600 ;
        RECT 196.600 21.800 197.500 22.200 ;
        RECT 197.100 21.100 197.500 21.800 ;
        RECT 201.400 21.100 201.800 24.800 ;
        RECT 202.200 24.800 203.300 25.100 ;
        RECT 202.200 21.100 202.600 24.800 ;
        RECT 0.600 15.700 1.000 19.900 ;
        RECT 2.800 18.200 3.200 19.900 ;
        RECT 2.200 17.900 3.200 18.200 ;
        RECT 5.000 17.900 5.400 19.900 ;
        RECT 7.100 17.900 7.700 19.900 ;
        RECT 2.200 17.500 2.600 17.900 ;
        RECT 5.000 17.600 5.300 17.900 ;
        RECT 3.900 17.300 5.700 17.600 ;
        RECT 7.000 17.500 7.400 17.900 ;
        RECT 3.900 17.200 4.300 17.300 ;
        RECT 5.300 17.200 5.700 17.300 ;
        RECT 2.200 16.500 2.600 16.600 ;
        RECT 4.500 16.500 4.900 16.600 ;
        RECT 2.200 16.200 4.900 16.500 ;
        RECT 5.200 16.500 6.300 16.800 ;
        RECT 5.200 15.900 5.500 16.500 ;
        RECT 5.900 16.400 6.300 16.500 ;
        RECT 7.100 16.600 7.800 17.000 ;
        RECT 7.100 16.100 7.400 16.600 ;
        RECT 3.100 15.700 5.500 15.900 ;
        RECT 0.600 15.600 5.500 15.700 ;
        RECT 6.200 15.800 7.400 16.100 ;
        RECT 0.600 15.500 3.500 15.600 ;
        RECT 0.600 15.400 3.400 15.500 ;
        RECT 6.200 15.200 6.500 15.800 ;
        RECT 9.400 15.600 9.800 19.900 ;
        RECT 10.200 16.200 10.600 19.900 ;
        RECT 11.800 16.200 12.200 19.900 ;
        RECT 10.200 15.900 12.200 16.200 ;
        RECT 12.600 15.900 13.000 19.900 ;
        RECT 13.700 16.300 14.100 19.900 ;
        RECT 13.700 15.900 14.600 16.300 ;
        RECT 7.700 15.300 9.800 15.600 ;
        RECT 7.700 15.200 8.100 15.300 ;
        RECT 3.800 15.100 4.200 15.200 ;
        RECT 5.400 15.100 5.800 15.200 ;
        RECT 1.700 14.800 5.800 15.100 ;
        RECT 6.200 14.800 6.600 15.200 ;
        RECT 8.500 14.900 8.900 15.000 ;
        RECT 1.700 14.700 2.100 14.800 ;
        RECT 2.500 14.200 2.900 14.300 ;
        RECT 6.200 14.200 6.500 14.800 ;
        RECT 7.000 14.600 8.900 14.900 ;
        RECT 7.000 14.500 7.400 14.600 ;
        RECT 1.000 13.900 6.500 14.200 ;
        RECT 9.400 14.100 9.800 15.300 ;
        RECT 10.600 15.200 11.000 15.400 ;
        RECT 12.600 15.200 12.900 15.900 ;
        RECT 10.200 14.900 11.000 15.200 ;
        RECT 11.800 14.900 13.000 15.200 ;
        RECT 10.200 14.800 10.600 14.900 ;
        RECT 10.200 14.100 10.600 14.200 ;
        RECT 1.000 13.800 1.800 13.900 ;
        RECT 0.600 11.100 1.000 13.500 ;
        RECT 3.100 12.800 3.400 13.900 ;
        RECT 5.900 13.800 6.300 13.900 ;
        RECT 9.400 13.800 10.600 14.100 ;
        RECT 11.000 13.800 11.400 14.600 ;
        RECT 9.400 13.600 9.800 13.800 ;
        RECT 7.900 13.300 9.800 13.600 ;
        RECT 7.900 13.200 8.300 13.300 ;
        RECT 2.200 12.100 2.600 12.500 ;
        RECT 3.000 12.400 3.400 12.800 ;
        RECT 3.900 12.700 4.300 12.800 ;
        RECT 3.900 12.400 5.300 12.700 ;
        RECT 5.000 12.100 5.300 12.400 ;
        RECT 7.000 12.100 7.400 12.500 ;
        RECT 2.200 11.800 3.200 12.100 ;
        RECT 2.800 11.100 3.200 11.800 ;
        RECT 5.000 11.100 5.400 12.100 ;
        RECT 7.000 11.800 7.700 12.100 ;
        RECT 7.100 11.100 7.700 11.800 ;
        RECT 9.400 11.100 9.800 13.300 ;
        RECT 11.800 13.200 12.100 14.900 ;
        RECT 12.600 14.800 13.000 14.900 ;
        RECT 13.400 14.800 13.800 15.600 ;
        RECT 14.200 14.200 14.500 15.900 ;
        RECT 15.800 15.700 16.200 19.900 ;
        RECT 18.000 18.200 18.400 19.900 ;
        RECT 17.400 17.900 18.400 18.200 ;
        RECT 20.200 17.900 20.600 19.900 ;
        RECT 22.300 17.900 22.900 19.900 ;
        RECT 17.400 17.500 17.800 17.900 ;
        RECT 20.200 17.600 20.500 17.900 ;
        RECT 19.100 17.300 20.900 17.600 ;
        RECT 22.200 17.500 22.600 17.900 ;
        RECT 19.100 17.200 19.500 17.300 ;
        RECT 20.500 17.200 20.900 17.300 ;
        RECT 17.400 16.500 17.800 16.600 ;
        RECT 19.700 16.500 20.100 16.600 ;
        RECT 17.400 16.200 20.100 16.500 ;
        RECT 20.400 16.500 21.500 16.800 ;
        RECT 20.400 15.900 20.700 16.500 ;
        RECT 21.100 16.400 21.500 16.500 ;
        RECT 22.300 16.600 23.000 17.000 ;
        RECT 22.300 16.100 22.600 16.600 ;
        RECT 18.300 15.700 20.700 15.900 ;
        RECT 15.800 15.600 20.700 15.700 ;
        RECT 21.400 15.800 22.600 16.100 ;
        RECT 15.800 15.500 18.700 15.600 ;
        RECT 15.800 15.400 18.600 15.500 ;
        RECT 19.000 15.100 19.400 15.200 ;
        RECT 16.900 14.800 19.400 15.100 ;
        RECT 20.600 15.100 21.000 15.200 ;
        RECT 21.400 15.100 21.700 15.800 ;
        RECT 24.600 15.600 25.000 19.900 ;
        RECT 26.700 16.200 27.100 19.900 ;
        RECT 27.400 16.800 27.800 17.200 ;
        RECT 27.500 16.200 27.800 16.800 ;
        RECT 26.700 15.900 27.200 16.200 ;
        RECT 27.500 15.900 28.200 16.200 ;
        RECT 22.900 15.300 25.000 15.600 ;
        RECT 22.900 15.200 23.300 15.300 ;
        RECT 20.600 14.800 21.700 15.100 ;
        RECT 23.700 14.900 24.100 15.000 ;
        RECT 16.900 14.700 17.300 14.800 ;
        RECT 17.700 14.200 18.100 14.300 ;
        RECT 21.400 14.200 21.700 14.800 ;
        RECT 22.200 14.600 24.100 14.900 ;
        RECT 22.200 14.500 22.600 14.600 ;
        RECT 14.200 13.800 14.600 14.200 ;
        RECT 16.200 13.900 21.700 14.200 ;
        RECT 16.200 13.800 17.000 13.900 ;
        RECT 11.800 11.100 12.200 13.200 ;
        RECT 12.600 13.100 13.000 13.200 ;
        RECT 14.200 13.100 14.500 13.800 ;
        RECT 12.600 12.800 14.500 13.100 ;
        RECT 12.500 12.400 12.900 12.800 ;
        RECT 14.200 12.100 14.500 12.800 ;
        RECT 15.000 12.400 15.400 13.200 ;
        RECT 14.200 11.100 14.600 12.100 ;
        RECT 15.800 11.100 16.200 13.500 ;
        RECT 18.300 12.800 18.600 13.900 ;
        RECT 21.100 13.800 21.500 13.900 ;
        RECT 24.600 13.600 25.000 15.300 ;
        RECT 26.900 15.200 27.200 15.900 ;
        RECT 27.800 15.800 28.200 15.900 ;
        RECT 28.600 15.800 29.000 16.600 ;
        RECT 26.200 14.400 26.600 15.200 ;
        RECT 26.900 14.800 27.400 15.200 ;
        RECT 27.800 15.100 28.100 15.800 ;
        RECT 29.400 15.100 29.800 19.900 ;
        RECT 32.300 16.200 32.700 19.900 ;
        RECT 33.000 16.800 33.400 17.200 ;
        RECT 33.100 16.200 33.400 16.800 ;
        RECT 32.300 15.900 32.800 16.200 ;
        RECT 33.100 15.900 33.800 16.200 ;
        RECT 27.800 14.800 29.800 15.100 ;
        RECT 26.900 14.200 27.200 14.800 ;
        RECT 25.400 14.100 25.800 14.200 ;
        RECT 25.400 13.800 26.200 14.100 ;
        RECT 26.900 13.800 28.200 14.200 ;
        RECT 25.800 13.600 26.200 13.800 ;
        RECT 23.100 13.300 25.000 13.600 ;
        RECT 23.100 13.200 23.500 13.300 ;
        RECT 17.400 12.100 17.800 12.500 ;
        RECT 18.200 12.400 18.600 12.800 ;
        RECT 19.100 12.700 19.500 12.800 ;
        RECT 19.100 12.400 20.500 12.700 ;
        RECT 20.200 12.100 20.500 12.400 ;
        RECT 22.200 12.100 22.600 12.500 ;
        RECT 17.400 11.800 18.400 12.100 ;
        RECT 18.000 11.100 18.400 11.800 ;
        RECT 20.200 11.100 20.600 12.100 ;
        RECT 22.200 11.800 22.900 12.100 ;
        RECT 22.300 11.100 22.900 11.800 ;
        RECT 24.600 11.100 25.000 13.300 ;
        RECT 25.500 13.100 27.300 13.300 ;
        RECT 27.800 13.100 28.100 13.800 ;
        RECT 29.400 13.100 29.800 14.800 ;
        RECT 31.800 14.400 32.200 15.200 ;
        RECT 32.500 14.200 32.800 15.900 ;
        RECT 33.400 15.800 33.800 15.900 ;
        RECT 34.200 15.800 34.600 16.600 ;
        RECT 33.400 15.100 33.700 15.800 ;
        RECT 35.000 15.100 35.400 19.900 ;
        RECT 33.400 14.800 35.400 15.100 ;
        RECT 30.200 13.400 30.600 14.200 ;
        RECT 31.000 14.100 31.400 14.200 ;
        RECT 31.000 13.800 31.800 14.100 ;
        RECT 32.500 13.800 33.800 14.200 ;
        RECT 31.400 13.600 31.800 13.800 ;
        RECT 31.100 13.100 32.900 13.300 ;
        RECT 33.400 13.100 33.700 13.800 ;
        RECT 35.000 13.100 35.400 14.800 ;
        RECT 35.800 13.400 36.200 14.200 ;
        RECT 25.400 13.000 27.400 13.100 ;
        RECT 25.400 11.100 25.800 13.000 ;
        RECT 27.000 11.100 27.400 13.000 ;
        RECT 27.800 11.100 28.200 13.100 ;
        RECT 28.900 12.800 29.800 13.100 ;
        RECT 31.000 13.000 33.000 13.100 ;
        RECT 28.900 11.100 29.300 12.800 ;
        RECT 31.000 11.100 31.400 13.000 ;
        RECT 32.600 11.100 33.000 13.000 ;
        RECT 33.400 11.100 33.800 13.100 ;
        RECT 34.500 12.800 35.400 13.100 ;
        RECT 34.500 11.100 34.900 12.800 ;
        RECT 36.600 12.400 37.000 13.200 ;
        RECT 37.400 11.100 37.800 19.900 ;
        RECT 38.200 14.800 38.600 15.200 ;
        RECT 38.200 14.200 38.500 14.800 ;
        RECT 38.200 13.400 38.600 14.200 ;
        RECT 39.000 13.100 39.400 19.900 ;
        RECT 39.800 15.800 40.200 16.600 ;
        RECT 40.600 15.700 41.000 19.900 ;
        RECT 42.800 18.200 43.200 19.900 ;
        RECT 42.200 17.900 43.200 18.200 ;
        RECT 45.000 17.900 45.400 19.900 ;
        RECT 47.100 17.900 47.700 19.900 ;
        RECT 42.200 17.500 42.600 17.900 ;
        RECT 45.000 17.600 45.300 17.900 ;
        RECT 43.900 17.300 45.700 17.600 ;
        RECT 47.000 17.500 47.400 17.900 ;
        RECT 43.900 17.200 44.300 17.300 ;
        RECT 45.300 17.200 45.700 17.300 ;
        RECT 42.200 16.500 42.600 16.600 ;
        RECT 44.500 16.500 44.900 16.600 ;
        RECT 42.200 16.200 44.900 16.500 ;
        RECT 45.200 16.500 46.300 16.800 ;
        RECT 45.200 15.900 45.500 16.500 ;
        RECT 45.900 16.400 46.300 16.500 ;
        RECT 47.100 16.600 47.800 17.000 ;
        RECT 47.100 16.100 47.400 16.600 ;
        RECT 43.100 15.700 45.500 15.900 ;
        RECT 40.600 15.600 45.500 15.700 ;
        RECT 46.200 15.800 47.400 16.100 ;
        RECT 40.600 15.500 43.500 15.600 ;
        RECT 40.600 15.400 43.400 15.500 ;
        RECT 43.800 15.100 44.200 15.200 ;
        RECT 41.700 14.800 44.200 15.100 ;
        RECT 41.700 14.700 42.100 14.800 ;
        RECT 42.500 14.200 42.900 14.300 ;
        RECT 46.200 14.200 46.500 15.800 ;
        RECT 49.400 15.600 49.800 19.900 ;
        RECT 53.100 16.200 53.500 19.900 ;
        RECT 53.800 16.800 54.200 17.200 ;
        RECT 53.900 16.200 54.200 16.800 ;
        RECT 53.100 15.900 53.600 16.200 ;
        RECT 53.900 15.900 54.600 16.200 ;
        RECT 47.700 15.300 49.800 15.600 ;
        RECT 47.700 15.200 48.100 15.300 ;
        RECT 48.500 14.900 48.900 15.000 ;
        RECT 47.000 14.600 48.900 14.900 ;
        RECT 47.000 14.500 47.400 14.600 ;
        RECT 41.000 13.900 46.500 14.200 ;
        RECT 41.000 13.800 41.800 13.900 ;
        RECT 39.000 12.800 39.900 13.100 ;
        RECT 39.500 12.200 39.900 12.800 ;
        RECT 39.500 11.800 40.200 12.200 ;
        RECT 39.500 11.100 39.900 11.800 ;
        RECT 40.600 11.100 41.000 13.500 ;
        RECT 43.100 12.800 43.400 13.900 ;
        RECT 43.800 13.800 44.200 13.900 ;
        RECT 45.900 13.800 46.300 13.900 ;
        RECT 49.400 13.600 49.800 15.300 ;
        RECT 53.300 15.200 53.600 15.900 ;
        RECT 54.200 15.800 54.600 15.900 ;
        RECT 55.000 15.800 55.400 16.600 ;
        RECT 52.600 14.400 53.000 15.200 ;
        RECT 53.300 14.800 53.800 15.200 ;
        RECT 54.200 15.100 54.500 15.800 ;
        RECT 55.800 15.100 56.200 19.900 ;
        RECT 58.700 19.200 59.100 19.900 ;
        RECT 58.700 18.800 59.400 19.200 ;
        RECT 58.700 16.300 59.100 18.800 ;
        RECT 58.200 15.900 59.100 16.300 ;
        RECT 60.100 16.300 60.500 19.900 ;
        RECT 60.100 15.900 61.000 16.300 ;
        RECT 54.200 14.800 56.200 15.100 ;
        RECT 53.300 14.200 53.600 14.800 ;
        RECT 51.800 14.100 52.200 14.200 ;
        RECT 51.800 13.800 52.600 14.100 ;
        RECT 53.300 13.800 54.600 14.200 ;
        RECT 52.200 13.600 52.600 13.800 ;
        RECT 47.900 13.300 49.800 13.600 ;
        RECT 47.900 13.200 48.300 13.300 ;
        RECT 42.200 12.100 42.600 12.500 ;
        RECT 43.000 12.400 43.400 12.800 ;
        RECT 43.900 12.700 44.300 12.800 ;
        RECT 43.900 12.400 45.300 12.700 ;
        RECT 45.000 12.100 45.300 12.400 ;
        RECT 47.000 12.100 47.400 12.500 ;
        RECT 42.200 11.800 43.200 12.100 ;
        RECT 42.800 11.100 43.200 11.800 ;
        RECT 45.000 11.100 45.400 12.100 ;
        RECT 47.000 11.800 47.700 12.100 ;
        RECT 47.100 11.100 47.700 11.800 ;
        RECT 49.400 11.100 49.800 13.300 ;
        RECT 51.900 13.100 53.700 13.300 ;
        RECT 54.200 13.100 54.500 13.800 ;
        RECT 55.800 13.100 56.200 14.800 ;
        RECT 58.300 14.200 58.600 15.900 ;
        RECT 59.000 15.100 59.400 15.600 ;
        RECT 59.800 15.100 60.200 15.600 ;
        RECT 59.000 14.800 60.200 15.100 ;
        RECT 60.600 15.100 60.900 15.900 ;
        RECT 62.200 15.600 62.600 19.900 ;
        RECT 64.300 17.900 64.900 19.900 ;
        RECT 66.600 17.900 67.000 19.900 ;
        RECT 68.800 18.200 69.200 19.900 ;
        RECT 68.800 17.900 69.800 18.200 ;
        RECT 64.600 17.500 65.000 17.900 ;
        RECT 66.700 17.600 67.000 17.900 ;
        RECT 66.300 17.300 68.100 17.600 ;
        RECT 69.400 17.500 69.800 17.900 ;
        RECT 66.300 17.200 66.700 17.300 ;
        RECT 67.700 17.200 68.100 17.300 ;
        RECT 64.200 16.600 64.900 17.000 ;
        RECT 64.600 16.100 64.900 16.600 ;
        RECT 65.700 16.500 66.800 16.800 ;
        RECT 65.700 16.400 66.100 16.500 ;
        RECT 64.600 15.800 65.800 16.100 ;
        RECT 62.200 15.300 64.300 15.600 ;
        RECT 60.600 14.800 61.700 15.100 ;
        RECT 56.600 13.400 57.000 14.200 ;
        RECT 58.200 13.800 58.600 14.200 ;
        RECT 51.800 13.000 53.800 13.100 ;
        RECT 51.800 11.100 52.200 13.000 ;
        RECT 53.400 11.100 53.800 13.000 ;
        RECT 54.200 11.100 54.600 13.100 ;
        RECT 55.300 12.800 56.200 13.100 ;
        RECT 55.300 11.100 55.700 12.800 ;
        RECT 57.400 12.400 57.800 13.200 ;
        RECT 58.300 12.100 58.600 13.800 ;
        RECT 58.200 11.100 58.600 12.100 ;
        RECT 60.600 14.200 60.900 14.800 ;
        RECT 61.400 14.200 61.700 14.800 ;
        RECT 60.600 13.800 61.000 14.200 ;
        RECT 61.400 13.800 61.800 14.200 ;
        RECT 60.600 12.100 60.900 13.800 ;
        RECT 62.200 13.600 62.600 15.300 ;
        RECT 63.900 15.200 64.300 15.300 ;
        RECT 63.100 14.900 63.500 15.000 ;
        RECT 63.100 14.600 65.000 14.900 ;
        RECT 64.600 14.500 65.000 14.600 ;
        RECT 65.500 14.200 65.800 15.800 ;
        RECT 66.500 15.900 66.800 16.500 ;
        RECT 67.100 16.500 67.500 16.600 ;
        RECT 69.400 16.500 69.800 16.600 ;
        RECT 67.100 16.200 69.800 16.500 ;
        RECT 66.500 15.700 68.900 15.900 ;
        RECT 71.000 15.700 71.400 19.900 ;
        RECT 73.100 16.200 73.500 19.900 ;
        RECT 73.800 16.800 74.200 17.200 ;
        RECT 73.900 16.200 74.200 16.800 ;
        RECT 76.300 16.200 76.700 19.900 ;
        RECT 77.000 16.800 77.400 17.200 ;
        RECT 77.100 16.200 77.400 16.800 ;
        RECT 73.100 15.900 73.600 16.200 ;
        RECT 73.900 15.900 74.600 16.200 ;
        RECT 76.300 15.900 76.800 16.200 ;
        RECT 77.100 15.900 77.800 16.200 ;
        RECT 79.500 15.900 80.500 19.900 ;
        RECT 66.500 15.600 71.400 15.700 ;
        RECT 68.500 15.500 71.400 15.600 ;
        RECT 68.600 15.400 71.400 15.500 ;
        RECT 67.800 15.100 68.200 15.200 ;
        RECT 67.800 14.800 70.300 15.100 ;
        RECT 68.600 14.700 69.000 14.800 ;
        RECT 69.900 14.700 70.300 14.800 ;
        RECT 72.600 14.400 73.000 15.200 ;
        RECT 69.100 14.200 69.500 14.300 ;
        RECT 73.300 14.200 73.600 15.900 ;
        RECT 74.200 15.800 74.600 15.900 ;
        RECT 75.800 14.400 76.200 15.200 ;
        RECT 76.500 14.200 76.800 15.900 ;
        RECT 77.400 15.800 77.800 15.900 ;
        RECT 65.500 13.900 71.000 14.200 ;
        RECT 65.700 13.800 66.100 13.900 ;
        RECT 62.200 13.300 64.100 13.600 ;
        RECT 61.400 12.400 61.800 13.200 ;
        RECT 60.600 11.100 61.000 12.100 ;
        RECT 62.200 11.100 62.600 13.300 ;
        RECT 63.700 13.200 64.100 13.300 ;
        RECT 68.600 12.800 68.900 13.900 ;
        RECT 70.200 13.800 71.000 13.900 ;
        RECT 71.800 14.100 72.200 14.200 ;
        RECT 71.800 13.800 72.600 14.100 ;
        RECT 73.300 13.800 74.600 14.200 ;
        RECT 75.000 14.100 75.400 14.200 ;
        RECT 76.500 14.100 77.800 14.200 ;
        RECT 78.200 14.100 78.600 14.600 ;
        RECT 79.000 14.400 79.400 15.200 ;
        RECT 79.900 14.200 80.200 15.900 ;
        RECT 80.600 15.100 81.000 15.200 ;
        RECT 81.400 15.100 81.800 15.200 ;
        RECT 80.600 14.800 81.800 15.100 ;
        RECT 80.600 14.400 81.000 14.800 ;
        RECT 79.800 14.100 80.200 14.200 ;
        RECT 81.400 14.100 81.800 14.200 ;
        RECT 75.000 13.800 75.800 14.100 ;
        RECT 76.500 13.800 78.600 14.100 ;
        RECT 79.000 13.800 80.200 14.100 ;
        RECT 81.000 13.800 81.800 14.100 ;
        RECT 72.200 13.600 72.600 13.800 ;
        RECT 67.700 12.700 68.100 12.800 ;
        RECT 64.600 12.100 65.000 12.500 ;
        RECT 66.700 12.400 68.100 12.700 ;
        RECT 68.600 12.400 69.000 12.800 ;
        RECT 66.700 12.100 67.000 12.400 ;
        RECT 69.400 12.100 69.800 12.500 ;
        RECT 64.300 11.800 65.000 12.100 ;
        RECT 64.300 11.100 64.900 11.800 ;
        RECT 66.600 11.100 67.000 12.100 ;
        RECT 68.800 11.800 69.800 12.100 ;
        RECT 68.800 11.100 69.200 11.800 ;
        RECT 71.000 11.100 71.400 13.500 ;
        RECT 71.900 13.100 73.700 13.300 ;
        RECT 74.200 13.100 74.500 13.800 ;
        RECT 75.400 13.600 75.800 13.800 ;
        RECT 75.100 13.100 76.900 13.300 ;
        RECT 77.400 13.100 77.700 13.800 ;
        RECT 79.000 13.100 79.300 13.800 ;
        RECT 81.000 13.600 81.400 13.800 ;
        RECT 79.900 13.100 81.700 13.300 ;
        RECT 71.800 13.000 73.800 13.100 ;
        RECT 71.800 11.100 72.200 13.000 ;
        RECT 73.400 11.100 73.800 13.000 ;
        RECT 74.200 11.100 74.600 13.100 ;
        RECT 75.000 13.000 77.000 13.100 ;
        RECT 75.000 11.100 75.400 13.000 ;
        RECT 76.600 11.100 77.000 13.000 ;
        RECT 77.400 11.100 77.800 13.100 ;
        RECT 78.200 11.400 78.600 13.100 ;
        RECT 79.000 11.700 79.400 13.100 ;
        RECT 79.800 13.000 81.800 13.100 ;
        RECT 79.800 11.400 80.200 13.000 ;
        RECT 78.200 11.100 80.200 11.400 ;
        RECT 81.400 11.100 81.800 13.000 ;
        RECT 82.200 12.400 82.600 13.200 ;
        RECT 83.000 11.100 83.400 19.900 ;
        RECT 84.600 15.100 85.000 19.900 ;
        RECT 86.600 16.800 87.000 17.200 ;
        RECT 85.400 15.800 85.800 16.600 ;
        RECT 86.600 16.200 86.900 16.800 ;
        RECT 87.300 16.200 87.700 19.900 ;
        RECT 86.200 15.900 86.900 16.200 ;
        RECT 87.200 15.900 87.700 16.200 ;
        RECT 86.200 15.800 86.600 15.900 ;
        RECT 86.200 15.100 86.500 15.800 ;
        RECT 84.600 14.800 86.500 15.100 ;
        RECT 83.800 13.400 84.200 14.200 ;
        RECT 84.600 13.100 85.000 14.800 ;
        RECT 87.200 14.200 87.500 15.900 ;
        RECT 89.400 15.700 89.800 19.900 ;
        RECT 91.600 18.200 92.000 19.900 ;
        RECT 91.000 17.900 92.000 18.200 ;
        RECT 93.800 17.900 94.200 19.900 ;
        RECT 95.900 17.900 96.500 19.900 ;
        RECT 91.000 17.500 91.400 17.900 ;
        RECT 93.800 17.600 94.100 17.900 ;
        RECT 92.700 17.300 94.500 17.600 ;
        RECT 95.800 17.500 96.200 17.900 ;
        RECT 92.700 17.200 93.100 17.300 ;
        RECT 94.100 17.200 94.500 17.300 ;
        RECT 91.000 16.500 91.400 16.600 ;
        RECT 93.300 16.500 93.700 16.600 ;
        RECT 91.000 16.200 93.700 16.500 ;
        RECT 94.000 16.500 95.100 16.800 ;
        RECT 94.000 15.900 94.300 16.500 ;
        RECT 94.700 16.400 95.100 16.500 ;
        RECT 95.900 16.600 96.600 17.000 ;
        RECT 95.900 16.100 96.200 16.600 ;
        RECT 91.900 15.700 94.300 15.900 ;
        RECT 89.400 15.600 94.300 15.700 ;
        RECT 95.000 15.800 96.200 16.100 ;
        RECT 89.400 15.500 92.300 15.600 ;
        RECT 89.400 15.400 92.200 15.500 ;
        RECT 87.800 14.400 88.200 15.200 ;
        RECT 92.600 15.100 93.000 15.200 ;
        RECT 94.200 15.100 94.600 15.200 ;
        RECT 90.500 14.800 94.600 15.100 ;
        RECT 90.500 14.700 90.900 14.800 ;
        RECT 91.300 14.200 91.700 14.300 ;
        RECT 95.000 14.200 95.300 15.800 ;
        RECT 98.200 15.600 98.600 19.900 ;
        RECT 96.500 15.300 98.600 15.600 ;
        RECT 96.500 15.200 96.900 15.300 ;
        RECT 97.300 14.900 97.700 15.000 ;
        RECT 95.800 14.600 97.700 14.900 ;
        RECT 95.800 14.500 96.200 14.600 ;
        RECT 86.200 13.800 87.500 14.200 ;
        RECT 88.600 14.100 89.000 14.200 ;
        RECT 88.200 13.800 89.000 14.100 ;
        RECT 89.800 13.900 95.300 14.200 ;
        RECT 89.800 13.800 90.600 13.900 ;
        RECT 86.300 13.100 86.600 13.800 ;
        RECT 88.200 13.600 88.600 13.800 ;
        RECT 87.100 13.100 88.900 13.300 ;
        RECT 84.600 12.800 85.500 13.100 ;
        RECT 85.100 11.100 85.500 12.800 ;
        RECT 86.200 11.100 86.600 13.100 ;
        RECT 87.000 13.000 89.000 13.100 ;
        RECT 87.000 11.100 87.400 13.000 ;
        RECT 88.600 11.100 89.000 13.000 ;
        RECT 89.400 11.100 89.800 13.500 ;
        RECT 91.900 13.200 92.200 13.900 ;
        RECT 94.700 13.800 95.100 13.900 ;
        RECT 98.200 13.600 98.600 15.300 ;
        RECT 96.700 13.300 98.600 13.600 ;
        RECT 96.700 13.200 97.100 13.300 ;
        RECT 91.000 12.100 91.400 12.500 ;
        RECT 91.800 12.400 92.200 13.200 ;
        RECT 92.700 12.700 93.100 12.800 ;
        RECT 92.700 12.400 94.100 12.700 ;
        RECT 93.800 12.100 94.100 12.400 ;
        RECT 95.800 12.100 96.200 12.500 ;
        RECT 91.000 11.800 92.000 12.100 ;
        RECT 91.600 11.100 92.000 11.800 ;
        RECT 93.800 11.100 94.200 12.100 ;
        RECT 95.800 11.800 96.500 12.100 ;
        RECT 95.900 11.100 96.500 11.800 ;
        RECT 98.200 11.100 98.600 13.300 ;
        RECT 99.000 11.100 99.400 19.900 ;
        RECT 101.900 16.300 102.300 19.900 ;
        RECT 101.400 15.900 102.300 16.300 ;
        RECT 101.500 15.100 101.800 15.900 ;
        RECT 104.600 15.600 105.000 19.900 ;
        RECT 106.700 17.900 107.300 19.900 ;
        RECT 109.000 17.900 109.400 19.900 ;
        RECT 111.200 18.200 111.600 19.900 ;
        RECT 111.200 17.900 112.200 18.200 ;
        RECT 107.000 17.500 107.400 17.900 ;
        RECT 109.100 17.600 109.400 17.900 ;
        RECT 108.700 17.300 110.500 17.600 ;
        RECT 111.800 17.500 112.200 17.900 ;
        RECT 108.700 17.200 109.100 17.300 ;
        RECT 110.100 17.200 110.500 17.300 ;
        RECT 106.600 16.600 107.300 17.000 ;
        RECT 107.000 16.100 107.300 16.600 ;
        RECT 108.100 16.500 109.200 16.800 ;
        RECT 108.100 16.400 108.500 16.500 ;
        RECT 107.000 15.800 108.200 16.100 ;
        RECT 99.800 14.800 101.800 15.100 ;
        RECT 102.200 14.800 102.600 15.600 ;
        RECT 104.600 15.300 106.700 15.600 ;
        RECT 99.800 14.200 100.100 14.800 ;
        RECT 101.500 14.200 101.800 14.800 ;
        RECT 99.800 13.800 100.200 14.200 ;
        RECT 101.400 13.800 101.800 14.200 ;
        RECT 99.800 12.400 100.200 13.200 ;
        RECT 100.600 12.400 101.000 13.200 ;
        RECT 101.500 12.100 101.800 13.800 ;
        RECT 101.400 11.100 101.800 12.100 ;
        RECT 104.600 13.600 105.000 15.300 ;
        RECT 106.300 15.200 106.700 15.300 ;
        RECT 105.500 14.900 105.900 15.000 ;
        RECT 105.500 14.600 107.400 14.900 ;
        RECT 107.000 14.500 107.400 14.600 ;
        RECT 107.900 14.200 108.200 15.800 ;
        RECT 108.900 15.900 109.200 16.500 ;
        RECT 109.500 16.500 109.900 16.600 ;
        RECT 111.800 16.500 112.200 16.600 ;
        RECT 109.500 16.200 112.200 16.500 ;
        RECT 108.900 15.700 111.300 15.900 ;
        RECT 113.400 15.700 113.800 19.900 ;
        RECT 108.900 15.600 113.800 15.700 ;
        RECT 110.900 15.500 113.800 15.600 ;
        RECT 111.000 15.400 113.800 15.500 ;
        RECT 110.200 15.100 110.600 15.200 ;
        RECT 115.000 15.100 115.400 19.900 ;
        RECT 117.000 16.800 117.400 17.200 ;
        RECT 115.800 15.800 116.200 16.600 ;
        RECT 117.000 16.200 117.300 16.800 ;
        RECT 117.700 16.200 118.100 19.900 ;
        RECT 116.600 15.900 117.300 16.200 ;
        RECT 117.600 15.900 118.100 16.200 ;
        RECT 116.600 15.800 117.000 15.900 ;
        RECT 116.600 15.100 116.900 15.800 ;
        RECT 117.600 15.200 117.900 15.900 ;
        RECT 119.800 15.700 120.200 19.900 ;
        RECT 122.000 18.200 122.400 19.900 ;
        RECT 121.400 17.900 122.400 18.200 ;
        RECT 124.200 17.900 124.600 19.900 ;
        RECT 126.300 17.900 126.900 19.900 ;
        RECT 121.400 17.500 121.800 17.900 ;
        RECT 124.200 17.600 124.500 17.900 ;
        RECT 123.100 17.300 124.900 17.600 ;
        RECT 126.200 17.500 126.600 17.900 ;
        RECT 123.100 17.200 123.500 17.300 ;
        RECT 124.500 17.200 124.900 17.300 ;
        RECT 121.400 16.500 121.800 16.600 ;
        RECT 123.700 16.500 124.100 16.600 ;
        RECT 121.400 16.200 124.100 16.500 ;
        RECT 124.400 16.500 125.500 16.800 ;
        RECT 124.400 15.900 124.700 16.500 ;
        RECT 125.100 16.400 125.500 16.500 ;
        RECT 126.300 16.600 127.000 17.000 ;
        RECT 126.300 16.100 126.600 16.600 ;
        RECT 122.300 15.700 124.700 15.900 ;
        RECT 119.800 15.600 124.700 15.700 ;
        RECT 125.400 15.800 126.600 16.100 ;
        RECT 119.800 15.500 122.700 15.600 ;
        RECT 119.800 15.400 122.600 15.500 ;
        RECT 110.200 14.800 112.700 15.100 ;
        RECT 112.300 14.700 112.700 14.800 ;
        RECT 115.000 14.800 116.900 15.100 ;
        RECT 117.400 14.800 117.900 15.200 ;
        RECT 111.500 14.200 111.900 14.300 ;
        RECT 107.900 13.900 113.400 14.200 ;
        RECT 108.100 13.800 108.500 13.900 ;
        RECT 110.200 13.800 110.600 13.900 ;
        RECT 104.600 13.300 106.500 13.600 ;
        RECT 104.600 11.100 105.000 13.300 ;
        RECT 106.100 13.200 106.500 13.300 ;
        RECT 111.000 12.800 111.300 13.900 ;
        RECT 112.600 13.800 113.400 13.900 ;
        RECT 110.100 12.700 110.500 12.800 ;
        RECT 107.000 12.100 107.400 12.500 ;
        RECT 109.100 12.400 110.500 12.700 ;
        RECT 111.000 12.400 111.400 12.800 ;
        RECT 109.100 12.100 109.400 12.400 ;
        RECT 111.800 12.100 112.200 12.500 ;
        RECT 106.700 11.800 107.400 12.100 ;
        RECT 106.700 11.100 107.300 11.800 ;
        RECT 109.000 11.100 109.400 12.100 ;
        RECT 111.200 11.800 112.200 12.100 ;
        RECT 111.200 11.100 111.600 11.800 ;
        RECT 113.400 11.100 113.800 13.500 ;
        RECT 114.200 13.400 114.600 14.200 ;
        RECT 115.000 13.100 115.400 14.800 ;
        RECT 117.600 14.200 117.900 14.800 ;
        RECT 118.200 14.400 118.600 15.200 ;
        RECT 123.000 15.100 123.400 15.200 ;
        RECT 120.900 14.800 123.400 15.100 ;
        RECT 120.900 14.700 121.300 14.800 ;
        RECT 122.200 14.700 122.600 14.800 ;
        RECT 121.700 14.200 122.100 14.300 ;
        RECT 125.400 14.200 125.700 15.800 ;
        RECT 128.600 15.600 129.000 19.900 ;
        RECT 130.200 15.600 130.600 19.900 ;
        RECT 131.800 15.600 132.200 19.900 ;
        RECT 133.400 15.600 133.800 19.900 ;
        RECT 135.000 15.600 135.400 19.900 ;
        RECT 126.900 15.300 129.000 15.600 ;
        RECT 126.900 15.200 127.300 15.300 ;
        RECT 127.700 14.900 128.100 15.000 ;
        RECT 126.200 14.600 128.100 14.900 ;
        RECT 126.200 14.500 126.600 14.600 ;
        RECT 116.600 13.800 117.900 14.200 ;
        RECT 119.000 14.100 119.400 14.200 ;
        RECT 118.600 13.800 119.400 14.100 ;
        RECT 120.200 13.900 125.700 14.200 ;
        RECT 120.200 13.800 121.000 13.900 ;
        RECT 116.700 13.100 117.000 13.800 ;
        RECT 118.600 13.600 119.000 13.800 ;
        RECT 117.500 13.100 119.300 13.300 ;
        RECT 115.000 12.800 115.900 13.100 ;
        RECT 115.500 11.100 115.900 12.800 ;
        RECT 116.600 11.100 117.000 13.100 ;
        RECT 117.400 13.000 119.400 13.100 ;
        RECT 117.400 11.100 117.800 13.000 ;
        RECT 119.000 11.100 119.400 13.000 ;
        RECT 119.800 11.100 120.200 13.500 ;
        RECT 122.300 12.800 122.600 13.900 ;
        RECT 125.100 13.800 125.500 13.900 ;
        RECT 128.600 13.600 129.000 15.300 ;
        RECT 127.000 13.300 129.000 13.600 ;
        RECT 129.400 15.200 130.600 15.600 ;
        RECT 131.100 15.200 132.200 15.600 ;
        RECT 132.700 15.200 133.800 15.600 ;
        RECT 134.500 15.200 135.400 15.600 ;
        RECT 136.600 17.500 137.000 19.500 ;
        RECT 136.600 15.800 136.900 17.500 ;
        RECT 138.700 16.400 139.100 19.900 ;
        RECT 138.700 16.100 139.500 16.400 ;
        RECT 142.700 16.300 143.100 19.900 ;
        RECT 136.600 15.500 138.500 15.800 ;
        RECT 129.400 13.800 129.800 15.200 ;
        RECT 131.100 14.500 131.500 15.200 ;
        RECT 132.700 14.500 133.100 15.200 ;
        RECT 134.500 14.500 134.900 15.200 ;
        RECT 130.200 14.100 131.500 14.500 ;
        RECT 131.900 14.100 133.100 14.500 ;
        RECT 133.600 14.100 134.900 14.500 ;
        RECT 136.600 14.400 137.000 15.200 ;
        RECT 137.400 14.400 137.800 15.200 ;
        RECT 138.200 14.500 138.500 15.500 ;
        RECT 131.100 13.800 131.500 14.100 ;
        RECT 132.700 13.800 133.100 14.100 ;
        RECT 134.500 13.800 134.900 14.100 ;
        RECT 138.200 14.100 138.900 14.500 ;
        RECT 139.200 14.200 139.500 16.100 ;
        RECT 142.200 15.900 143.100 16.300 ;
        RECT 143.800 15.900 144.200 19.900 ;
        RECT 144.600 16.200 145.000 19.900 ;
        RECT 146.200 16.200 146.600 19.900 ;
        RECT 144.600 15.900 146.600 16.200 ;
        RECT 139.800 15.100 140.200 15.600 ;
        RECT 141.400 15.100 141.800 15.200 ;
        RECT 139.800 14.800 141.800 15.100 ;
        RECT 142.300 14.200 142.600 15.900 ;
        RECT 143.000 14.800 143.400 15.600 ;
        RECT 143.900 15.200 144.200 15.900 ;
        RECT 147.000 15.600 147.400 19.900 ;
        RECT 149.100 17.900 149.700 19.900 ;
        RECT 151.400 17.900 151.800 19.900 ;
        RECT 153.600 18.200 154.000 19.900 ;
        RECT 153.600 17.900 154.600 18.200 ;
        RECT 149.400 17.500 149.800 17.900 ;
        RECT 151.500 17.600 151.800 17.900 ;
        RECT 151.100 17.300 152.900 17.600 ;
        RECT 154.200 17.500 154.600 17.900 ;
        RECT 151.100 17.200 151.500 17.300 ;
        RECT 152.500 17.200 152.900 17.300 ;
        RECT 148.600 17.000 149.300 17.200 ;
        RECT 148.600 16.800 149.700 17.000 ;
        RECT 149.000 16.600 149.700 16.800 ;
        RECT 149.400 16.100 149.700 16.600 ;
        RECT 150.500 16.500 151.600 16.800 ;
        RECT 150.500 16.400 150.900 16.500 ;
        RECT 149.400 15.800 150.600 16.100 ;
        RECT 145.800 15.200 146.200 15.400 ;
        RECT 147.000 15.300 149.100 15.600 ;
        RECT 143.800 14.900 145.000 15.200 ;
        RECT 145.800 14.900 146.600 15.200 ;
        RECT 143.800 14.800 144.200 14.900 ;
        RECT 138.200 13.900 138.700 14.100 ;
        RECT 129.400 13.400 130.600 13.800 ;
        RECT 131.100 13.400 132.200 13.800 ;
        RECT 132.700 13.400 133.800 13.800 ;
        RECT 134.500 13.400 135.400 13.800 ;
        RECT 127.000 13.200 127.500 13.300 ;
        RECT 125.400 13.100 125.800 13.200 ;
        RECT 127.000 13.100 127.400 13.200 ;
        RECT 125.400 12.800 127.400 13.100 ;
        RECT 121.400 12.100 121.800 12.500 ;
        RECT 122.200 12.400 122.600 12.800 ;
        RECT 123.100 12.700 123.500 12.800 ;
        RECT 123.100 12.400 124.500 12.700 ;
        RECT 124.200 12.100 124.500 12.400 ;
        RECT 126.200 12.100 126.600 12.500 ;
        RECT 121.400 11.800 122.400 12.100 ;
        RECT 122.000 11.100 122.400 11.800 ;
        RECT 124.200 11.100 124.600 12.100 ;
        RECT 126.200 11.800 126.900 12.100 ;
        RECT 126.300 11.100 126.900 11.800 ;
        RECT 128.600 11.100 129.000 13.300 ;
        RECT 130.200 11.100 130.600 13.400 ;
        RECT 131.800 11.100 132.200 13.400 ;
        RECT 133.400 11.100 133.800 13.400 ;
        RECT 135.000 11.100 135.400 13.400 ;
        RECT 136.600 13.600 138.700 13.900 ;
        RECT 139.200 13.800 140.200 14.200 ;
        RECT 142.200 13.800 142.600 14.200 ;
        RECT 136.600 12.500 136.900 13.600 ;
        RECT 139.200 13.500 139.500 13.800 ;
        RECT 139.100 13.300 139.500 13.500 ;
        RECT 138.700 13.000 139.500 13.300 ;
        RECT 136.600 11.500 137.000 12.500 ;
        RECT 138.700 12.200 139.100 13.000 ;
        RECT 141.400 12.400 141.800 13.200 ;
        RECT 142.300 13.100 142.600 13.800 ;
        RECT 144.700 13.200 145.000 14.900 ;
        RECT 146.200 14.800 146.600 14.900 ;
        RECT 145.400 13.800 145.800 14.600 ;
        RECT 143.800 13.100 144.200 13.200 ;
        RECT 142.200 12.800 144.200 13.100 ;
        RECT 138.700 11.800 139.400 12.200 ;
        RECT 142.300 12.100 142.600 12.800 ;
        RECT 143.900 12.400 144.300 12.800 ;
        RECT 138.700 11.500 139.100 11.800 ;
        RECT 142.200 11.100 142.600 12.100 ;
        RECT 144.600 11.100 145.000 13.200 ;
        RECT 147.000 13.600 147.400 15.300 ;
        RECT 148.700 15.200 149.100 15.300 ;
        RECT 150.300 15.200 150.600 15.800 ;
        RECT 151.300 15.900 151.600 16.500 ;
        RECT 151.900 16.500 152.300 16.600 ;
        RECT 154.200 16.500 154.600 16.600 ;
        RECT 151.900 16.200 154.600 16.500 ;
        RECT 151.300 15.700 153.700 15.900 ;
        RECT 155.800 15.700 156.200 19.900 ;
        RECT 159.500 16.300 159.900 19.900 ;
        RECT 159.000 15.900 159.900 16.300 ;
        RECT 160.600 15.900 161.000 19.900 ;
        RECT 161.400 16.200 161.800 19.900 ;
        RECT 163.000 16.200 163.400 19.900 ;
        RECT 165.100 16.300 165.500 19.900 ;
        RECT 161.400 15.900 163.400 16.200 ;
        RECT 164.600 15.900 165.500 16.300 ;
        RECT 166.200 15.900 166.600 19.900 ;
        RECT 167.000 16.200 167.400 19.900 ;
        RECT 168.600 16.200 169.000 19.900 ;
        RECT 167.000 15.900 169.000 16.200 ;
        RECT 151.300 15.600 156.200 15.700 ;
        RECT 153.300 15.500 156.200 15.600 ;
        RECT 153.400 15.400 156.200 15.500 ;
        RECT 147.900 14.900 148.300 15.000 ;
        RECT 147.900 14.600 149.800 14.900 ;
        RECT 150.200 14.800 150.600 15.200 ;
        RECT 151.000 15.100 151.400 15.200 ;
        RECT 152.600 15.100 153.000 15.200 ;
        RECT 151.000 14.800 155.100 15.100 ;
        RECT 149.400 14.500 149.800 14.600 ;
        RECT 150.300 14.200 150.600 14.800 ;
        RECT 154.700 14.700 155.100 14.800 ;
        RECT 153.900 14.200 154.300 14.300 ;
        RECT 159.100 14.200 159.400 15.900 ;
        RECT 159.800 14.800 160.200 15.600 ;
        RECT 160.700 15.200 161.000 15.900 ;
        RECT 162.600 15.200 163.000 15.400 ;
        RECT 160.600 14.900 161.800 15.200 ;
        RECT 162.600 14.900 163.400 15.200 ;
        RECT 160.600 14.800 161.000 14.900 ;
        RECT 150.300 13.900 155.800 14.200 ;
        RECT 150.500 13.800 150.900 13.900 ;
        RECT 147.000 13.300 148.900 13.600 ;
        RECT 147.000 11.100 147.400 13.300 ;
        RECT 148.500 13.200 148.900 13.300 ;
        RECT 153.400 12.800 153.700 13.900 ;
        RECT 155.000 13.800 155.800 13.900 ;
        RECT 159.000 13.800 159.400 14.200 ;
        RECT 152.500 12.700 152.900 12.800 ;
        RECT 149.400 12.100 149.800 12.500 ;
        RECT 151.500 12.400 152.900 12.700 ;
        RECT 153.400 12.400 153.800 12.800 ;
        RECT 151.500 12.100 151.800 12.400 ;
        RECT 154.200 12.100 154.600 12.500 ;
        RECT 149.100 11.800 149.800 12.100 ;
        RECT 149.100 11.100 149.700 11.800 ;
        RECT 151.400 11.100 151.800 12.100 ;
        RECT 153.600 11.800 154.600 12.100 ;
        RECT 153.600 11.100 154.000 11.800 ;
        RECT 155.800 11.100 156.200 13.500 ;
        RECT 156.600 13.100 157.000 13.200 ;
        RECT 158.200 13.100 158.600 13.200 ;
        RECT 159.100 13.100 159.400 13.800 ;
        RECT 160.600 13.100 161.000 13.200 ;
        RECT 161.500 13.100 161.800 14.900 ;
        RECT 163.000 14.800 163.400 14.900 ;
        RECT 162.200 13.800 162.600 14.600 ;
        RECT 164.700 14.200 165.000 15.900 ;
        RECT 165.400 14.800 165.800 15.600 ;
        RECT 166.300 15.200 166.600 15.900 ;
        RECT 170.200 15.600 170.600 19.900 ;
        RECT 171.800 15.600 172.200 19.900 ;
        RECT 173.400 15.600 173.800 19.900 ;
        RECT 175.000 15.600 175.400 19.900 ;
        RECT 177.900 16.300 178.300 19.900 ;
        RECT 177.400 15.900 178.300 16.300 ;
        RECT 179.000 15.900 179.400 19.900 ;
        RECT 179.800 16.200 180.200 19.900 ;
        RECT 181.400 16.200 181.800 19.900 ;
        RECT 183.500 16.300 183.900 19.900 ;
        RECT 179.800 15.900 181.800 16.200 ;
        RECT 183.000 15.900 183.900 16.300 ;
        RECT 184.600 15.900 185.000 19.900 ;
        RECT 185.400 16.200 185.800 19.900 ;
        RECT 187.000 16.200 187.400 19.900 ;
        RECT 185.400 15.900 187.400 16.200 ;
        RECT 168.200 15.200 168.600 15.400 ;
        RECT 170.200 15.200 171.100 15.600 ;
        RECT 171.800 15.200 172.900 15.600 ;
        RECT 173.400 15.200 174.500 15.600 ;
        RECT 175.000 15.200 176.200 15.600 ;
        RECT 166.200 14.900 167.400 15.200 ;
        RECT 168.200 14.900 169.000 15.200 ;
        RECT 166.200 14.800 166.600 14.900 ;
        RECT 164.600 13.800 165.000 14.200 ;
        RECT 156.600 12.800 158.600 13.100 ;
        RECT 159.000 12.800 161.000 13.100 ;
        RECT 158.200 12.400 158.600 12.800 ;
        RECT 159.100 12.100 159.400 12.800 ;
        RECT 160.700 12.400 161.100 12.800 ;
        RECT 159.000 11.100 159.400 12.100 ;
        RECT 161.400 11.100 161.800 13.100 ;
        RECT 163.800 12.400 164.200 13.200 ;
        RECT 164.700 13.100 165.000 13.800 ;
        RECT 166.200 13.100 166.600 13.200 ;
        RECT 167.100 13.100 167.400 14.900 ;
        RECT 168.600 14.800 169.000 14.900 ;
        RECT 167.800 13.800 168.200 14.600 ;
        RECT 170.700 14.500 171.100 15.200 ;
        RECT 172.500 14.500 172.900 15.200 ;
        RECT 174.100 14.500 174.500 15.200 ;
        RECT 170.700 14.100 172.000 14.500 ;
        RECT 172.500 14.100 173.700 14.500 ;
        RECT 174.100 14.100 175.400 14.500 ;
        RECT 170.700 13.800 171.100 14.100 ;
        RECT 172.500 13.800 172.900 14.100 ;
        RECT 174.100 13.800 174.500 14.100 ;
        RECT 175.800 13.800 176.200 15.200 ;
        RECT 177.500 14.200 177.800 15.900 ;
        RECT 178.200 14.800 178.600 15.600 ;
        RECT 179.100 15.200 179.400 15.900 ;
        RECT 181.000 15.200 181.400 15.400 ;
        RECT 179.000 14.900 180.200 15.200 ;
        RECT 181.000 14.900 181.800 15.200 ;
        RECT 179.000 14.800 179.400 14.900 ;
        RECT 177.400 13.800 177.800 14.200 ;
        RECT 164.600 12.800 166.600 13.100 ;
        RECT 164.700 12.100 165.000 12.800 ;
        RECT 166.300 12.400 166.700 12.800 ;
        RECT 164.600 11.100 165.000 12.100 ;
        RECT 167.000 11.100 167.400 13.100 ;
        RECT 170.200 13.400 171.100 13.800 ;
        RECT 171.800 13.400 172.900 13.800 ;
        RECT 173.400 13.400 174.500 13.800 ;
        RECT 175.000 13.400 176.200 13.800 ;
        RECT 170.200 11.100 170.600 13.400 ;
        RECT 171.800 11.100 172.200 13.400 ;
        RECT 173.400 11.100 173.800 13.400 ;
        RECT 175.000 11.100 175.400 13.400 ;
        RECT 176.600 12.400 177.000 13.200 ;
        RECT 177.500 13.100 177.800 13.800 ;
        RECT 179.000 13.100 179.400 13.200 ;
        RECT 179.900 13.100 180.200 14.900 ;
        RECT 181.400 14.800 181.800 14.900 ;
        RECT 180.600 13.800 181.000 14.600 ;
        RECT 183.100 14.200 183.400 15.900 ;
        RECT 183.800 14.800 184.200 15.600 ;
        RECT 184.700 15.200 185.000 15.900 ;
        RECT 187.800 15.700 188.200 19.900 ;
        RECT 190.000 18.200 190.400 19.900 ;
        RECT 189.400 17.900 190.400 18.200 ;
        RECT 192.200 17.900 192.600 19.900 ;
        RECT 194.300 17.900 194.900 19.900 ;
        RECT 189.400 17.500 189.800 17.900 ;
        RECT 192.200 17.600 192.500 17.900 ;
        RECT 191.100 17.300 192.900 17.600 ;
        RECT 194.200 17.500 194.600 17.900 ;
        RECT 191.100 17.200 191.500 17.300 ;
        RECT 192.500 17.200 192.900 17.300 ;
        RECT 189.400 16.500 189.800 16.600 ;
        RECT 191.700 16.500 192.100 16.600 ;
        RECT 189.400 16.200 192.100 16.500 ;
        RECT 192.400 16.500 193.500 16.800 ;
        RECT 192.400 15.900 192.700 16.500 ;
        RECT 193.100 16.400 193.500 16.500 ;
        RECT 194.300 16.600 195.000 17.000 ;
        RECT 194.300 16.100 194.600 16.600 ;
        RECT 190.300 15.700 192.700 15.900 ;
        RECT 187.800 15.600 192.700 15.700 ;
        RECT 193.400 15.800 194.600 16.100 ;
        RECT 187.800 15.500 190.700 15.600 ;
        RECT 187.800 15.400 190.600 15.500 ;
        RECT 186.600 15.200 187.000 15.400 ;
        RECT 184.600 14.900 185.800 15.200 ;
        RECT 186.600 14.900 187.400 15.200 ;
        RECT 191.000 15.100 191.400 15.200 ;
        RECT 184.600 14.800 185.000 14.900 ;
        RECT 183.000 13.800 183.400 14.200 ;
        RECT 177.400 12.800 179.400 13.100 ;
        RECT 177.500 12.100 177.800 12.800 ;
        RECT 179.100 12.400 179.500 12.800 ;
        RECT 177.400 11.100 177.800 12.100 ;
        RECT 179.800 11.100 180.200 13.100 ;
        RECT 182.200 12.400 182.600 13.200 ;
        RECT 183.100 13.100 183.400 13.800 ;
        RECT 184.600 13.100 185.000 13.200 ;
        RECT 185.500 13.100 185.800 14.900 ;
        RECT 187.000 14.800 187.400 14.900 ;
        RECT 188.900 14.800 191.400 15.100 ;
        RECT 188.900 14.700 189.300 14.800 ;
        RECT 190.200 14.700 190.600 14.800 ;
        RECT 186.200 13.800 186.600 14.600 ;
        RECT 189.700 14.200 190.100 14.300 ;
        RECT 193.400 14.200 193.700 15.800 ;
        RECT 196.600 15.600 197.000 19.900 ;
        RECT 197.400 16.200 197.800 19.900 ;
        RECT 197.400 15.900 198.500 16.200 ;
        RECT 194.900 15.300 197.000 15.600 ;
        RECT 194.900 15.200 195.300 15.300 ;
        RECT 195.700 14.900 196.100 15.000 ;
        RECT 194.200 14.600 196.100 14.900 ;
        RECT 194.200 14.500 194.600 14.600 ;
        RECT 188.200 13.900 193.700 14.200 ;
        RECT 188.200 13.800 189.000 13.900 ;
        RECT 183.000 12.800 185.000 13.100 ;
        RECT 183.100 12.100 183.400 12.800 ;
        RECT 184.700 12.400 185.100 12.800 ;
        RECT 183.000 11.100 183.400 12.100 ;
        RECT 185.400 11.100 185.800 13.100 ;
        RECT 187.800 11.100 188.200 13.500 ;
        RECT 190.300 12.800 190.600 13.900 ;
        RECT 193.100 13.800 193.500 13.900 ;
        RECT 196.600 13.600 197.000 15.300 ;
        RECT 198.200 15.600 198.500 15.900 ;
        RECT 198.200 15.200 198.800 15.600 ;
        RECT 197.400 14.400 197.800 15.200 ;
        RECT 198.200 13.700 198.500 15.200 ;
        RECT 195.100 13.300 197.000 13.600 ;
        RECT 195.100 13.200 195.500 13.300 ;
        RECT 189.400 12.100 189.800 12.500 ;
        RECT 190.200 12.400 190.600 12.800 ;
        RECT 191.100 12.700 191.500 12.800 ;
        RECT 191.100 12.400 192.500 12.700 ;
        RECT 192.200 12.100 192.500 12.400 ;
        RECT 194.200 12.100 194.600 12.500 ;
        RECT 189.400 11.800 190.400 12.100 ;
        RECT 190.000 11.100 190.400 11.800 ;
        RECT 192.200 11.100 192.600 12.100 ;
        RECT 194.200 11.800 194.900 12.100 ;
        RECT 194.300 11.100 194.900 11.800 ;
        RECT 196.600 11.100 197.000 13.300 ;
        RECT 197.400 13.400 198.500 13.700 ;
        RECT 197.400 11.100 197.800 13.400 ;
        RECT 199.800 11.100 200.200 19.900 ;
        RECT 201.400 16.200 201.800 19.900 ;
        RECT 201.400 15.900 202.500 16.200 ;
        RECT 202.200 15.600 202.500 15.900 ;
        RECT 202.200 15.200 202.800 15.600 ;
        RECT 200.600 15.100 201.000 15.200 ;
        RECT 201.400 15.100 201.800 15.200 ;
        RECT 200.600 14.800 201.800 15.100 ;
        RECT 201.400 14.400 201.800 14.800 ;
        RECT 202.200 13.700 202.500 15.200 ;
        RECT 201.400 13.400 202.500 13.700 ;
        RECT 200.600 12.400 201.000 13.200 ;
        RECT 201.400 11.100 201.800 13.400 ;
        RECT 1.400 7.600 1.800 9.900 ;
        RECT 3.000 7.600 3.400 9.900 ;
        RECT 4.600 7.600 5.000 9.900 ;
        RECT 6.200 7.600 6.600 9.900 ;
        RECT 8.600 7.600 9.000 9.900 ;
        RECT 10.200 7.600 10.600 9.900 ;
        RECT 11.800 7.600 12.200 9.900 ;
        RECT 13.400 7.600 13.800 9.900 ;
        RECT 1.400 7.200 2.300 7.600 ;
        RECT 3.000 7.200 4.100 7.600 ;
        RECT 4.600 7.200 5.700 7.600 ;
        RECT 6.200 7.200 7.400 7.600 ;
        RECT 8.600 7.200 9.500 7.600 ;
        RECT 10.200 7.200 11.300 7.600 ;
        RECT 11.800 7.200 12.900 7.600 ;
        RECT 13.400 7.200 14.600 7.600 ;
        RECT 15.000 7.500 15.400 9.900 ;
        RECT 17.200 9.200 17.600 9.900 ;
        RECT 16.600 8.900 17.600 9.200 ;
        RECT 19.400 8.900 19.800 9.900 ;
        RECT 21.500 9.200 22.100 9.900 ;
        RECT 21.400 8.900 22.100 9.200 ;
        RECT 16.600 8.500 17.000 8.900 ;
        RECT 19.400 8.600 19.700 8.900 ;
        RECT 17.400 8.200 17.800 8.600 ;
        RECT 18.300 8.300 19.700 8.600 ;
        RECT 21.400 8.500 21.800 8.900 ;
        RECT 18.300 8.200 18.700 8.300 ;
        RECT 1.900 6.900 2.300 7.200 ;
        RECT 3.700 6.900 4.100 7.200 ;
        RECT 5.300 6.900 5.700 7.200 ;
        RECT 1.900 6.500 3.200 6.900 ;
        RECT 3.700 6.500 4.900 6.900 ;
        RECT 5.300 6.500 6.600 6.900 ;
        RECT 1.900 5.800 2.300 6.500 ;
        RECT 3.700 5.800 4.100 6.500 ;
        RECT 5.300 5.800 5.700 6.500 ;
        RECT 7.000 5.800 7.400 7.200 ;
        RECT 9.100 6.900 9.500 7.200 ;
        RECT 10.900 6.900 11.300 7.200 ;
        RECT 12.500 6.900 12.900 7.200 ;
        RECT 9.100 6.500 10.400 6.900 ;
        RECT 10.900 6.500 12.100 6.900 ;
        RECT 12.500 6.500 13.800 6.900 ;
        RECT 9.100 5.800 9.500 6.500 ;
        RECT 10.900 5.800 11.300 6.500 ;
        RECT 12.500 5.800 12.900 6.500 ;
        RECT 14.200 5.800 14.600 7.200 ;
        RECT 15.400 7.100 16.200 7.200 ;
        RECT 17.500 7.100 17.800 8.200 ;
        RECT 23.800 8.100 24.200 9.900 ;
        RECT 25.400 8.900 25.800 9.900 ;
        RECT 24.600 8.100 25.000 8.600 ;
        RECT 25.500 8.100 25.800 8.900 ;
        RECT 27.100 8.200 27.500 8.600 ;
        RECT 27.000 8.100 27.400 8.200 ;
        RECT 23.800 7.800 25.000 8.100 ;
        RECT 25.400 7.800 27.400 8.100 ;
        RECT 27.800 7.900 28.200 9.900 ;
        RECT 22.300 7.700 22.700 7.800 ;
        RECT 23.800 7.700 24.200 7.800 ;
        RECT 22.300 7.400 24.200 7.700 ;
        RECT 20.300 7.100 20.700 7.200 ;
        RECT 15.400 6.800 20.900 7.100 ;
        RECT 16.900 6.700 17.300 6.800 ;
        RECT 16.100 6.200 16.500 6.300 ;
        RECT 16.100 5.900 18.600 6.200 ;
        RECT 18.200 5.800 18.600 5.900 ;
        RECT 1.400 5.400 2.300 5.800 ;
        RECT 3.000 5.400 4.100 5.800 ;
        RECT 4.600 5.400 5.700 5.800 ;
        RECT 6.200 5.400 7.400 5.800 ;
        RECT 8.600 5.400 9.500 5.800 ;
        RECT 10.200 5.400 11.300 5.800 ;
        RECT 11.800 5.400 12.900 5.800 ;
        RECT 13.400 5.400 14.600 5.800 ;
        RECT 15.000 5.500 17.800 5.600 ;
        RECT 15.000 5.400 17.900 5.500 ;
        RECT 1.400 1.100 1.800 5.400 ;
        RECT 3.000 1.100 3.400 5.400 ;
        RECT 4.600 1.100 5.000 5.400 ;
        RECT 6.200 1.100 6.600 5.400 ;
        RECT 8.600 1.100 9.000 5.400 ;
        RECT 10.200 1.100 10.600 5.400 ;
        RECT 11.800 1.100 12.200 5.400 ;
        RECT 13.400 1.100 13.800 5.400 ;
        RECT 15.000 5.300 19.900 5.400 ;
        RECT 15.000 1.100 15.400 5.300 ;
        RECT 17.500 5.100 19.900 5.300 ;
        RECT 16.600 4.500 19.300 4.800 ;
        RECT 16.600 4.400 17.000 4.500 ;
        RECT 18.900 4.400 19.300 4.500 ;
        RECT 19.600 4.500 19.900 5.100 ;
        RECT 20.600 5.200 20.900 6.800 ;
        RECT 21.400 6.400 21.800 6.500 ;
        RECT 21.400 6.100 23.300 6.400 ;
        RECT 22.900 6.000 23.300 6.100 ;
        RECT 22.100 5.700 22.500 5.800 ;
        RECT 23.800 5.700 24.200 7.400 ;
        RECT 25.500 7.200 25.800 7.800 ;
        RECT 25.400 6.800 25.800 7.200 ;
        RECT 22.100 5.400 24.200 5.700 ;
        RECT 20.600 4.900 21.800 5.200 ;
        RECT 20.300 4.500 20.700 4.600 ;
        RECT 19.600 4.200 20.700 4.500 ;
        RECT 21.500 4.400 21.800 4.900 ;
        RECT 21.500 4.000 22.200 4.400 ;
        RECT 18.300 3.700 18.700 3.800 ;
        RECT 19.700 3.700 20.100 3.800 ;
        RECT 16.600 3.100 17.000 3.500 ;
        RECT 18.300 3.400 20.100 3.700 ;
        RECT 19.400 3.100 19.700 3.400 ;
        RECT 21.400 3.100 21.800 3.500 ;
        RECT 16.600 2.800 17.600 3.100 ;
        RECT 17.200 1.100 17.600 2.800 ;
        RECT 19.400 1.100 19.800 3.100 ;
        RECT 21.500 1.100 22.100 3.100 ;
        RECT 23.800 1.100 24.200 5.400 ;
        RECT 25.500 5.100 25.800 6.800 ;
        RECT 27.000 6.800 27.400 7.200 ;
        RECT 27.000 6.200 27.300 6.800 ;
        RECT 26.200 5.400 26.600 6.200 ;
        RECT 27.000 6.100 27.400 6.200 ;
        RECT 27.900 6.100 28.200 7.900 ;
        RECT 30.200 7.500 30.600 9.900 ;
        RECT 32.400 9.200 32.800 9.900 ;
        RECT 31.800 8.900 32.800 9.200 ;
        RECT 34.600 8.900 35.000 9.900 ;
        RECT 36.700 9.200 37.300 9.900 ;
        RECT 36.600 8.900 37.300 9.200 ;
        RECT 31.800 8.500 32.200 8.900 ;
        RECT 34.600 8.600 34.900 8.900 ;
        RECT 32.600 8.200 33.000 8.600 ;
        RECT 33.500 8.300 34.900 8.600 ;
        RECT 36.600 8.500 37.000 8.900 ;
        RECT 33.500 8.200 33.900 8.300 ;
        RECT 28.600 6.400 29.000 7.200 ;
        RECT 30.600 7.100 31.400 7.200 ;
        RECT 32.700 7.100 33.000 8.200 ;
        RECT 37.500 7.700 37.900 7.800 ;
        RECT 39.000 7.700 39.400 9.900 ;
        RECT 39.800 7.900 40.200 9.900 ;
        RECT 40.600 8.000 41.000 9.900 ;
        RECT 42.200 8.000 42.600 9.900 ;
        RECT 40.600 7.900 42.600 8.000 ;
        RECT 37.500 7.400 39.400 7.700 ;
        RECT 35.500 7.100 35.900 7.200 ;
        RECT 30.600 6.800 36.100 7.100 ;
        RECT 32.100 6.700 32.500 6.800 ;
        RECT 31.300 6.200 31.700 6.300 ;
        RECT 29.400 6.100 29.800 6.200 ;
        RECT 27.000 5.800 28.200 6.100 ;
        RECT 29.000 5.800 29.800 6.100 ;
        RECT 31.300 5.900 33.800 6.200 ;
        RECT 33.400 5.800 33.800 5.900 ;
        RECT 27.100 5.100 27.400 5.800 ;
        RECT 29.000 5.600 29.400 5.800 ;
        RECT 30.200 5.500 33.000 5.600 ;
        RECT 30.200 5.400 33.100 5.500 ;
        RECT 30.200 5.300 35.100 5.400 ;
        RECT 25.400 4.700 26.300 5.100 ;
        RECT 25.900 1.100 26.300 4.700 ;
        RECT 27.000 1.100 27.400 5.100 ;
        RECT 27.800 4.800 29.800 5.100 ;
        RECT 27.800 1.100 28.200 4.800 ;
        RECT 29.400 1.100 29.800 4.800 ;
        RECT 30.200 1.100 30.600 5.300 ;
        RECT 32.700 5.100 35.100 5.300 ;
        RECT 31.800 4.500 34.500 4.800 ;
        RECT 31.800 4.400 32.200 4.500 ;
        RECT 34.100 4.400 34.500 4.500 ;
        RECT 34.800 4.500 35.100 5.100 ;
        RECT 35.800 5.200 36.100 6.800 ;
        RECT 36.600 6.400 37.000 6.500 ;
        RECT 36.600 6.100 38.500 6.400 ;
        RECT 38.100 6.000 38.500 6.100 ;
        RECT 37.300 5.700 37.700 5.800 ;
        RECT 39.000 5.700 39.400 7.400 ;
        RECT 39.900 7.200 40.200 7.900 ;
        RECT 40.700 7.700 42.500 7.900 ;
        RECT 43.000 7.700 43.400 9.900 ;
        RECT 45.100 9.200 45.700 9.900 ;
        RECT 45.100 8.900 45.800 9.200 ;
        RECT 47.400 8.900 47.800 9.900 ;
        RECT 49.600 9.200 50.000 9.900 ;
        RECT 49.600 8.900 50.600 9.200 ;
        RECT 45.400 8.500 45.800 8.900 ;
        RECT 47.500 8.600 47.800 8.900 ;
        RECT 47.500 8.300 48.900 8.600 ;
        RECT 48.500 8.200 48.900 8.300 ;
        RECT 49.400 8.200 49.800 8.600 ;
        RECT 50.200 8.500 50.600 8.900 ;
        RECT 44.500 7.700 44.900 7.800 ;
        RECT 43.000 7.400 44.900 7.700 ;
        RECT 41.800 7.200 42.200 7.400 ;
        RECT 39.800 6.800 41.100 7.200 ;
        RECT 41.800 6.900 42.600 7.200 ;
        RECT 42.200 6.800 42.600 6.900 ;
        RECT 37.300 5.400 39.400 5.700 ;
        RECT 35.800 4.900 37.000 5.200 ;
        RECT 35.500 4.500 35.900 4.600 ;
        RECT 34.800 4.200 35.900 4.500 ;
        RECT 36.700 4.400 37.000 4.900 ;
        RECT 36.700 4.000 37.400 4.400 ;
        RECT 33.500 3.700 33.900 3.800 ;
        RECT 34.900 3.700 35.300 3.800 ;
        RECT 31.800 3.100 32.200 3.500 ;
        RECT 33.500 3.400 35.300 3.700 ;
        RECT 34.600 3.100 34.900 3.400 ;
        RECT 36.600 3.100 37.000 3.500 ;
        RECT 31.800 2.800 32.800 3.100 ;
        RECT 32.400 1.100 32.800 2.800 ;
        RECT 34.600 1.100 35.000 3.100 ;
        RECT 36.700 1.100 37.300 3.100 ;
        RECT 39.000 1.100 39.400 5.400 ;
        RECT 40.800 5.200 41.100 6.800 ;
        RECT 41.400 5.800 41.800 6.600 ;
        RECT 43.000 5.700 43.400 7.400 ;
        RECT 46.500 7.100 46.900 7.200 ;
        RECT 49.400 7.100 49.700 8.200 ;
        RECT 51.800 7.500 52.200 9.900 ;
        RECT 54.200 7.500 54.600 9.900 ;
        RECT 56.400 9.200 56.800 9.900 ;
        RECT 55.800 8.900 56.800 9.200 ;
        RECT 58.600 8.900 59.000 9.900 ;
        RECT 60.700 9.200 61.300 9.900 ;
        RECT 60.600 8.900 61.300 9.200 ;
        RECT 55.800 8.500 56.200 8.900 ;
        RECT 58.600 8.600 58.900 8.900 ;
        RECT 56.600 8.200 57.000 8.600 ;
        RECT 57.500 8.300 58.900 8.600 ;
        RECT 60.600 8.500 61.000 8.900 ;
        RECT 57.500 8.200 57.900 8.300 ;
        RECT 51.000 7.100 51.800 7.200 ;
        RECT 54.600 7.100 55.400 7.200 ;
        RECT 56.700 7.100 57.000 8.200 ;
        RECT 59.800 7.800 60.200 8.200 ;
        RECT 61.400 7.800 61.800 8.200 ;
        RECT 59.800 7.200 60.100 7.800 ;
        RECT 61.400 7.700 61.900 7.800 ;
        RECT 63.000 7.700 63.400 9.900 ;
        RECT 65.100 8.200 65.500 9.900 ;
        RECT 61.400 7.400 63.400 7.700 ;
        RECT 64.600 7.900 65.500 8.200 ;
        RECT 66.200 7.900 66.600 9.900 ;
        RECT 67.000 8.000 67.400 9.900 ;
        RECT 68.600 8.000 69.000 9.900 ;
        RECT 67.000 7.900 69.000 8.000 ;
        RECT 59.500 7.100 60.100 7.200 ;
        RECT 46.300 6.800 60.100 7.100 ;
        RECT 45.400 6.400 45.800 6.500 ;
        RECT 43.900 6.100 45.800 6.400 ;
        RECT 46.300 6.200 46.600 6.800 ;
        RECT 49.900 6.700 50.300 6.800 ;
        RECT 56.100 6.700 56.500 6.800 ;
        RECT 50.700 6.200 51.100 6.300 ;
        RECT 43.900 6.000 44.300 6.100 ;
        RECT 46.200 5.800 46.600 6.200 ;
        RECT 48.600 5.900 51.100 6.200 ;
        RECT 55.300 6.200 55.700 6.300 ;
        RECT 55.300 5.900 57.800 6.200 ;
        RECT 48.600 5.800 49.000 5.900 ;
        RECT 57.400 5.800 57.800 5.900 ;
        RECT 44.700 5.700 45.100 5.800 ;
        RECT 43.000 5.400 45.100 5.700 ;
        RECT 39.800 5.100 40.200 5.200 ;
        RECT 39.800 4.800 40.500 5.100 ;
        RECT 40.800 4.800 41.800 5.200 ;
        RECT 40.200 4.200 40.500 4.800 ;
        RECT 40.200 3.800 40.600 4.200 ;
        RECT 40.900 1.100 41.300 4.800 ;
        RECT 43.000 1.100 43.400 5.400 ;
        RECT 46.300 5.200 46.600 5.800 ;
        RECT 49.400 5.500 52.200 5.600 ;
        RECT 49.300 5.400 52.200 5.500 ;
        RECT 45.400 4.900 46.600 5.200 ;
        RECT 47.300 5.300 52.200 5.400 ;
        RECT 47.300 5.100 49.700 5.300 ;
        RECT 45.400 4.400 45.700 4.900 ;
        RECT 45.000 4.000 45.700 4.400 ;
        RECT 46.500 4.500 46.900 4.600 ;
        RECT 47.300 4.500 47.600 5.100 ;
        RECT 46.500 4.200 47.600 4.500 ;
        RECT 47.900 4.500 50.600 4.800 ;
        RECT 47.900 4.400 48.300 4.500 ;
        RECT 50.200 4.400 50.600 4.500 ;
        RECT 47.100 3.700 47.500 3.800 ;
        RECT 48.500 3.700 48.900 3.800 ;
        RECT 45.400 3.100 45.800 3.500 ;
        RECT 47.100 3.400 48.900 3.700 ;
        RECT 47.500 3.100 47.800 3.400 ;
        RECT 50.200 3.100 50.600 3.500 ;
        RECT 45.100 1.100 45.700 3.100 ;
        RECT 47.400 1.100 47.800 3.100 ;
        RECT 49.600 2.800 50.600 3.100 ;
        RECT 49.600 1.100 50.000 2.800 ;
        RECT 51.800 1.100 52.200 5.300 ;
        RECT 54.200 5.500 57.000 5.600 ;
        RECT 54.200 5.400 57.100 5.500 ;
        RECT 54.200 5.300 59.100 5.400 ;
        RECT 54.200 1.100 54.600 5.300 ;
        RECT 56.700 5.100 59.100 5.300 ;
        RECT 55.800 4.500 58.500 4.800 ;
        RECT 55.800 4.400 56.200 4.500 ;
        RECT 58.100 4.400 58.500 4.500 ;
        RECT 58.800 4.500 59.100 5.100 ;
        RECT 59.800 5.200 60.100 6.800 ;
        RECT 63.000 7.100 63.400 7.400 ;
        RECT 63.800 7.100 64.200 7.600 ;
        RECT 63.000 6.800 64.200 7.100 ;
        RECT 60.600 6.400 61.000 6.500 ;
        RECT 60.600 6.100 62.500 6.400 ;
        RECT 62.100 6.000 62.500 6.100 ;
        RECT 61.300 5.700 61.700 5.800 ;
        RECT 63.000 5.700 63.400 6.800 ;
        RECT 61.300 5.400 63.400 5.700 ;
        RECT 59.800 4.900 61.000 5.200 ;
        RECT 59.500 4.500 59.900 4.600 ;
        RECT 58.800 4.200 59.900 4.500 ;
        RECT 60.700 4.400 61.000 4.900 ;
        RECT 60.700 4.000 61.400 4.400 ;
        RECT 57.500 3.700 57.900 3.800 ;
        RECT 58.900 3.700 59.300 3.800 ;
        RECT 55.800 3.100 56.200 3.500 ;
        RECT 57.500 3.400 59.300 3.700 ;
        RECT 58.600 3.100 58.900 3.400 ;
        RECT 60.600 3.100 61.000 3.500 ;
        RECT 55.800 2.800 56.800 3.100 ;
        RECT 56.400 1.100 56.800 2.800 ;
        RECT 58.600 1.100 59.000 3.100 ;
        RECT 60.700 1.100 61.300 3.100 ;
        RECT 63.000 1.100 63.400 5.400 ;
        RECT 64.600 6.100 65.000 7.900 ;
        RECT 66.300 7.200 66.600 7.900 ;
        RECT 67.100 7.700 68.900 7.900 ;
        RECT 69.400 7.500 69.800 9.900 ;
        RECT 71.600 9.200 72.000 9.900 ;
        RECT 71.000 8.900 72.000 9.200 ;
        RECT 73.800 8.900 74.200 9.900 ;
        RECT 75.900 9.200 76.500 9.900 ;
        RECT 75.800 8.900 76.500 9.200 ;
        RECT 71.000 8.500 71.400 8.900 ;
        RECT 73.800 8.600 74.100 8.900 ;
        RECT 71.800 8.200 72.200 8.600 ;
        RECT 72.700 8.300 74.100 8.600 ;
        RECT 75.800 8.500 76.200 8.900 ;
        RECT 72.700 8.200 73.100 8.300 ;
        RECT 68.200 7.200 68.600 7.400 ;
        RECT 65.400 7.100 65.800 7.200 ;
        RECT 66.200 7.100 67.500 7.200 ;
        RECT 65.400 6.800 67.500 7.100 ;
        RECT 68.200 6.900 69.000 7.200 ;
        RECT 68.600 6.800 69.000 6.900 ;
        RECT 69.800 7.100 70.600 7.200 ;
        RECT 71.900 7.100 72.200 8.200 ;
        RECT 76.700 7.700 77.100 7.800 ;
        RECT 78.200 7.700 78.600 9.900 ;
        RECT 79.300 9.200 79.700 9.900 ;
        RECT 79.000 8.800 79.700 9.200 ;
        RECT 79.300 8.200 79.700 8.800 ;
        RECT 79.300 7.900 80.200 8.200 ;
        RECT 76.700 7.400 78.600 7.700 ;
        RECT 74.700 7.100 75.100 7.200 ;
        RECT 69.800 6.800 75.300 7.100 ;
        RECT 64.600 5.800 66.500 6.100 ;
        RECT 64.600 1.100 65.000 5.800 ;
        RECT 66.200 5.200 66.500 5.800 ;
        RECT 65.400 4.400 65.800 5.200 ;
        RECT 66.200 5.100 66.600 5.200 ;
        RECT 67.200 5.100 67.500 6.800 ;
        RECT 71.300 6.700 71.700 6.800 ;
        RECT 67.800 5.800 68.200 6.600 ;
        RECT 70.500 6.200 70.900 6.300 ;
        RECT 70.500 6.100 73.000 6.200 ;
        RECT 74.200 6.100 74.600 6.200 ;
        RECT 70.500 5.900 74.600 6.100 ;
        RECT 72.600 5.800 74.600 5.900 ;
        RECT 69.400 5.500 72.200 5.600 ;
        RECT 69.400 5.400 72.300 5.500 ;
        RECT 69.400 5.300 74.300 5.400 ;
        RECT 66.200 4.800 66.900 5.100 ;
        RECT 67.200 4.800 67.700 5.100 ;
        RECT 66.600 4.200 66.900 4.800 ;
        RECT 66.600 3.800 67.000 4.200 ;
        RECT 67.300 1.100 67.700 4.800 ;
        RECT 69.400 1.100 69.800 5.300 ;
        RECT 71.900 5.100 74.300 5.300 ;
        RECT 71.000 4.500 73.700 4.800 ;
        RECT 71.000 4.400 71.400 4.500 ;
        RECT 73.300 4.400 73.700 4.500 ;
        RECT 74.000 4.500 74.300 5.100 ;
        RECT 75.000 5.200 75.300 6.800 ;
        RECT 75.800 6.400 76.200 6.500 ;
        RECT 75.800 6.100 77.700 6.400 ;
        RECT 77.300 6.000 77.700 6.100 ;
        RECT 76.500 5.700 76.900 5.800 ;
        RECT 78.200 5.700 78.600 7.400 ;
        RECT 76.500 5.400 78.600 5.700 ;
        RECT 75.000 4.900 76.200 5.200 ;
        RECT 74.700 4.500 75.100 4.600 ;
        RECT 74.000 4.200 75.100 4.500 ;
        RECT 75.900 4.400 76.200 4.900 ;
        RECT 75.900 4.000 76.600 4.400 ;
        RECT 72.700 3.700 73.100 3.800 ;
        RECT 74.100 3.700 74.500 3.800 ;
        RECT 71.000 3.100 71.400 3.500 ;
        RECT 72.700 3.400 74.500 3.700 ;
        RECT 73.800 3.100 74.100 3.400 ;
        RECT 75.800 3.100 76.200 3.500 ;
        RECT 71.000 2.800 72.000 3.100 ;
        RECT 71.600 1.100 72.000 2.800 ;
        RECT 73.800 1.100 74.200 3.100 ;
        RECT 75.900 1.100 76.500 3.100 ;
        RECT 78.200 1.100 78.600 5.400 ;
        RECT 79.000 4.400 79.400 5.200 ;
        RECT 79.800 1.100 80.200 7.900 ;
        RECT 81.400 7.700 81.800 9.900 ;
        RECT 83.500 9.200 84.100 9.900 ;
        RECT 83.500 8.900 84.200 9.200 ;
        RECT 85.800 8.900 86.200 9.900 ;
        RECT 88.000 9.200 88.400 9.900 ;
        RECT 88.000 8.900 89.000 9.200 ;
        RECT 83.800 8.500 84.200 8.900 ;
        RECT 85.900 8.600 86.200 8.900 ;
        RECT 85.900 8.300 87.300 8.600 ;
        RECT 86.900 8.200 87.300 8.300 ;
        RECT 87.800 8.200 88.200 8.600 ;
        RECT 88.600 8.500 89.000 8.900 ;
        RECT 82.900 7.700 83.300 7.800 ;
        RECT 80.600 6.800 81.000 7.600 ;
        RECT 81.400 7.400 83.300 7.700 ;
        RECT 81.400 5.700 81.800 7.400 ;
        RECT 82.200 6.800 82.600 7.400 ;
        RECT 84.900 7.100 85.300 7.200 ;
        RECT 87.800 7.100 88.100 8.200 ;
        RECT 90.200 7.500 90.600 9.900 ;
        RECT 91.000 7.700 91.400 9.900 ;
        RECT 93.100 9.200 93.700 9.900 ;
        RECT 93.100 8.900 93.800 9.200 ;
        RECT 95.400 8.900 95.800 9.900 ;
        RECT 97.600 9.200 98.000 9.900 ;
        RECT 97.600 8.900 98.600 9.200 ;
        RECT 93.400 8.500 93.800 8.900 ;
        RECT 95.500 8.600 95.800 8.900 ;
        RECT 95.500 8.300 96.900 8.600 ;
        RECT 96.500 8.200 96.900 8.300 ;
        RECT 97.400 8.200 97.800 8.600 ;
        RECT 98.200 8.500 98.600 8.900 ;
        RECT 92.500 7.700 92.900 7.800 ;
        RECT 91.000 7.400 92.900 7.700 ;
        RECT 89.400 7.100 90.200 7.200 ;
        RECT 84.700 6.800 90.200 7.100 ;
        RECT 83.800 6.400 84.200 6.500 ;
        RECT 82.300 6.100 84.200 6.400 ;
        RECT 84.700 6.200 85.000 6.800 ;
        RECT 88.300 6.700 88.700 6.800 ;
        RECT 89.100 6.200 89.500 6.300 ;
        RECT 82.300 6.000 82.700 6.100 ;
        RECT 84.600 5.800 85.000 6.200 ;
        RECT 87.000 5.900 89.500 6.200 ;
        RECT 87.000 5.800 87.400 5.900 ;
        RECT 83.100 5.700 83.500 5.800 ;
        RECT 81.400 5.400 83.500 5.700 ;
        RECT 81.400 1.100 81.800 5.400 ;
        RECT 84.700 5.200 85.000 5.800 ;
        RECT 91.000 5.700 91.400 7.400 ;
        RECT 94.500 7.100 94.900 7.200 ;
        RECT 97.400 7.100 97.700 8.200 ;
        RECT 99.800 7.500 100.200 9.900 ;
        RECT 102.200 7.700 102.600 9.900 ;
        RECT 104.300 9.200 104.900 9.900 ;
        RECT 104.300 8.900 105.000 9.200 ;
        RECT 106.600 8.900 107.000 9.900 ;
        RECT 108.800 9.200 109.200 9.900 ;
        RECT 108.800 8.900 109.800 9.200 ;
        RECT 104.600 8.500 105.000 8.900 ;
        RECT 106.700 8.600 107.000 8.900 ;
        RECT 106.700 8.300 108.100 8.600 ;
        RECT 107.700 8.200 108.100 8.300 ;
        RECT 108.600 8.200 109.000 8.600 ;
        RECT 109.400 8.500 109.800 8.900 ;
        RECT 103.700 7.700 104.100 7.800 ;
        RECT 102.200 7.400 104.100 7.700 ;
        RECT 99.000 7.100 99.800 7.200 ;
        RECT 94.300 6.800 99.800 7.100 ;
        RECT 93.400 6.400 93.800 6.500 ;
        RECT 91.900 6.100 93.800 6.400 ;
        RECT 94.300 6.200 94.600 6.800 ;
        RECT 97.900 6.700 98.300 6.800 ;
        RECT 98.700 6.200 99.100 6.300 ;
        RECT 91.900 6.000 92.300 6.100 ;
        RECT 94.200 5.800 94.600 6.200 ;
        RECT 96.600 5.900 99.100 6.200 ;
        RECT 96.600 5.800 97.000 5.900 ;
        RECT 92.700 5.700 93.100 5.800 ;
        RECT 87.800 5.500 90.600 5.600 ;
        RECT 87.700 5.400 90.600 5.500 ;
        RECT 83.800 4.900 85.000 5.200 ;
        RECT 85.700 5.300 90.600 5.400 ;
        RECT 85.700 5.100 88.100 5.300 ;
        RECT 83.800 4.400 84.100 4.900 ;
        RECT 83.400 4.000 84.100 4.400 ;
        RECT 84.900 4.500 85.300 4.600 ;
        RECT 85.700 4.500 86.000 5.100 ;
        RECT 84.900 4.200 86.000 4.500 ;
        RECT 86.300 4.500 89.000 4.800 ;
        RECT 86.300 4.400 86.700 4.500 ;
        RECT 88.600 4.400 89.000 4.500 ;
        RECT 85.500 3.700 85.900 3.800 ;
        RECT 86.900 3.700 87.300 3.800 ;
        RECT 83.800 3.100 84.200 3.500 ;
        RECT 85.500 3.400 87.300 3.700 ;
        RECT 85.900 3.100 86.200 3.400 ;
        RECT 88.600 3.100 89.000 3.500 ;
        RECT 83.500 1.100 84.100 3.100 ;
        RECT 85.800 1.100 86.200 3.100 ;
        RECT 88.000 2.800 89.000 3.100 ;
        RECT 88.000 1.100 88.400 2.800 ;
        RECT 90.200 1.100 90.600 5.300 ;
        RECT 91.000 5.400 93.100 5.700 ;
        RECT 91.000 1.100 91.400 5.400 ;
        RECT 94.300 5.200 94.600 5.800 ;
        RECT 102.200 5.700 102.600 7.400 ;
        RECT 105.700 7.100 106.100 7.200 ;
        RECT 108.600 7.100 108.900 8.200 ;
        RECT 111.000 7.500 111.400 9.900 ;
        RECT 113.100 8.200 113.500 9.900 ;
        RECT 112.600 7.900 113.500 8.200 ;
        RECT 114.200 7.900 114.600 9.900 ;
        RECT 115.000 8.000 115.400 9.900 ;
        RECT 116.600 8.000 117.000 9.900 ;
        RECT 115.000 7.900 117.000 8.000 ;
        RECT 118.200 8.900 118.600 9.900 ;
        RECT 110.200 7.100 111.000 7.200 ;
        RECT 105.500 6.800 111.000 7.100 ;
        RECT 111.800 6.800 112.200 7.600 ;
        RECT 104.600 6.400 105.000 6.500 ;
        RECT 103.100 6.100 105.000 6.400 ;
        RECT 105.500 6.200 105.800 6.800 ;
        RECT 109.100 6.700 109.500 6.800 ;
        RECT 108.600 6.200 109.000 6.300 ;
        RECT 109.900 6.200 110.300 6.300 ;
        RECT 103.100 6.000 103.500 6.100 ;
        RECT 105.400 5.800 105.800 6.200 ;
        RECT 107.800 5.900 110.300 6.200 ;
        RECT 112.600 6.100 113.000 7.900 ;
        RECT 114.300 7.200 114.600 7.900 ;
        RECT 115.100 7.700 116.900 7.900 ;
        RECT 116.200 7.200 116.600 7.400 ;
        RECT 118.200 7.200 118.500 8.900 ;
        RECT 119.000 7.800 119.400 8.600 ;
        RECT 119.900 8.200 120.300 8.600 ;
        RECT 119.800 7.800 120.200 8.200 ;
        RECT 120.600 7.900 121.000 9.900 ;
        RECT 113.400 7.100 113.800 7.200 ;
        RECT 114.200 7.100 115.500 7.200 ;
        RECT 113.400 6.800 115.500 7.100 ;
        RECT 116.200 6.900 117.000 7.200 ;
        RECT 116.600 6.800 117.000 6.900 ;
        RECT 118.200 7.100 118.600 7.200 ;
        RECT 119.800 7.100 120.100 7.800 ;
        RECT 118.200 6.800 120.100 7.100 ;
        RECT 107.800 5.800 108.200 5.900 ;
        RECT 112.600 5.800 114.500 6.100 ;
        RECT 103.900 5.700 104.300 5.800 ;
        RECT 97.400 5.500 100.200 5.600 ;
        RECT 97.300 5.400 100.200 5.500 ;
        RECT 93.400 4.900 94.600 5.200 ;
        RECT 95.300 5.300 100.200 5.400 ;
        RECT 95.300 5.100 97.700 5.300 ;
        RECT 93.400 4.400 93.700 4.900 ;
        RECT 93.000 4.000 93.700 4.400 ;
        RECT 94.500 4.500 94.900 4.600 ;
        RECT 95.300 4.500 95.600 5.100 ;
        RECT 94.500 4.200 95.600 4.500 ;
        RECT 95.900 4.500 98.600 4.800 ;
        RECT 95.900 4.400 96.300 4.500 ;
        RECT 98.200 4.400 98.600 4.500 ;
        RECT 95.100 3.700 95.500 3.800 ;
        RECT 96.500 3.700 96.900 3.800 ;
        RECT 93.400 3.100 93.800 3.500 ;
        RECT 95.100 3.400 96.900 3.700 ;
        RECT 95.500 3.100 95.800 3.400 ;
        RECT 98.200 3.100 98.600 3.500 ;
        RECT 93.100 1.100 93.700 3.100 ;
        RECT 95.400 1.100 95.800 3.100 ;
        RECT 97.600 2.800 98.600 3.100 ;
        RECT 97.600 1.100 98.000 2.800 ;
        RECT 99.800 1.100 100.200 5.300 ;
        RECT 102.200 5.400 104.300 5.700 ;
        RECT 102.200 1.100 102.600 5.400 ;
        RECT 105.500 5.200 105.800 5.800 ;
        RECT 108.600 5.500 111.400 5.600 ;
        RECT 108.500 5.400 111.400 5.500 ;
        RECT 104.600 4.900 105.800 5.200 ;
        RECT 106.500 5.300 111.400 5.400 ;
        RECT 106.500 5.100 108.900 5.300 ;
        RECT 104.600 4.400 104.900 4.900 ;
        RECT 104.200 4.000 104.900 4.400 ;
        RECT 105.700 4.500 106.100 4.600 ;
        RECT 106.500 4.500 106.800 5.100 ;
        RECT 105.700 4.200 106.800 4.500 ;
        RECT 107.100 4.500 109.800 4.800 ;
        RECT 107.100 4.400 107.500 4.500 ;
        RECT 109.400 4.400 109.800 4.500 ;
        RECT 106.300 3.700 106.700 3.800 ;
        RECT 107.700 3.700 108.100 3.800 ;
        RECT 104.600 3.100 105.000 3.500 ;
        RECT 106.300 3.400 108.100 3.700 ;
        RECT 106.700 3.100 107.000 3.400 ;
        RECT 109.400 3.100 109.800 3.500 ;
        RECT 104.300 1.100 104.900 3.100 ;
        RECT 106.600 1.100 107.000 3.100 ;
        RECT 108.800 2.800 109.800 3.100 ;
        RECT 108.800 1.100 109.200 2.800 ;
        RECT 111.000 1.100 111.400 5.300 ;
        RECT 112.600 1.100 113.000 5.800 ;
        RECT 114.200 5.200 114.500 5.800 ;
        RECT 113.400 4.400 113.800 5.200 ;
        RECT 114.200 5.100 114.600 5.200 ;
        RECT 115.200 5.100 115.500 6.800 ;
        RECT 115.800 5.800 116.200 6.600 ;
        RECT 117.400 5.400 117.800 6.200 ;
        RECT 118.200 5.100 118.500 6.800 ;
        RECT 120.700 6.200 121.000 7.900 ;
        RECT 123.000 7.700 123.400 9.900 ;
        RECT 125.100 9.200 125.700 9.900 ;
        RECT 125.100 8.900 125.800 9.200 ;
        RECT 127.400 8.900 127.800 9.900 ;
        RECT 129.600 9.200 130.000 9.900 ;
        RECT 129.600 8.900 130.600 9.200 ;
        RECT 125.400 8.500 125.800 8.900 ;
        RECT 127.500 8.600 127.800 8.900 ;
        RECT 127.500 8.300 128.900 8.600 ;
        RECT 128.500 8.200 128.900 8.300 ;
        RECT 129.400 8.200 129.800 8.600 ;
        RECT 130.200 8.500 130.600 8.900 ;
        RECT 124.500 7.700 124.900 7.800 ;
        RECT 123.000 7.400 124.900 7.700 ;
        RECT 121.400 6.400 121.800 7.200 ;
        RECT 119.800 6.100 120.200 6.200 ;
        RECT 120.600 6.100 121.000 6.200 ;
        RECT 122.200 6.100 122.600 6.200 ;
        RECT 119.800 5.800 121.000 6.100 ;
        RECT 121.800 5.800 122.600 6.100 ;
        RECT 119.900 5.100 120.200 5.800 ;
        RECT 121.800 5.600 122.200 5.800 ;
        RECT 123.000 5.700 123.400 7.400 ;
        RECT 126.500 7.100 126.900 7.200 ;
        RECT 129.400 7.100 129.700 8.200 ;
        RECT 131.800 7.500 132.200 9.900 ;
        RECT 131.000 7.100 131.800 7.200 ;
        RECT 126.300 6.800 131.800 7.100 ;
        RECT 125.400 6.400 125.800 6.500 ;
        RECT 123.900 6.100 125.800 6.400 ;
        RECT 123.900 6.000 124.300 6.100 ;
        RECT 124.700 5.700 125.100 5.800 ;
        RECT 123.000 5.400 125.100 5.700 ;
        RECT 114.200 4.800 114.900 5.100 ;
        RECT 115.200 4.800 115.700 5.100 ;
        RECT 114.600 4.200 114.900 4.800 ;
        RECT 114.600 3.800 115.000 4.200 ;
        RECT 115.300 1.100 115.700 4.800 ;
        RECT 117.700 4.700 118.600 5.100 ;
        RECT 117.700 1.100 118.100 4.700 ;
        RECT 119.800 1.100 120.200 5.100 ;
        RECT 120.600 4.800 122.600 5.100 ;
        RECT 120.600 1.100 121.000 4.800 ;
        RECT 122.200 1.100 122.600 4.800 ;
        RECT 123.000 1.100 123.400 5.400 ;
        RECT 126.300 5.200 126.600 6.800 ;
        RECT 129.900 6.700 130.300 6.800 ;
        RECT 130.700 6.200 131.100 6.300 ;
        RECT 127.000 6.100 127.400 6.200 ;
        RECT 128.600 6.100 131.100 6.200 ;
        RECT 127.000 5.900 131.100 6.100 ;
        RECT 127.000 5.800 129.000 5.900 ;
        RECT 129.400 5.500 132.200 5.600 ;
        RECT 129.300 5.400 132.200 5.500 ;
        RECT 125.400 4.900 126.600 5.200 ;
        RECT 127.300 5.300 132.200 5.400 ;
        RECT 127.300 5.100 129.700 5.300 ;
        RECT 125.400 4.400 125.700 4.900 ;
        RECT 125.000 4.000 125.700 4.400 ;
        RECT 126.500 4.500 126.900 4.600 ;
        RECT 127.300 4.500 127.600 5.100 ;
        RECT 126.500 4.200 127.600 4.500 ;
        RECT 127.900 4.500 130.600 4.800 ;
        RECT 127.900 4.400 128.300 4.500 ;
        RECT 130.200 4.400 130.600 4.500 ;
        RECT 127.100 3.700 127.500 3.800 ;
        RECT 128.500 3.700 128.900 3.800 ;
        RECT 125.400 3.100 125.800 3.500 ;
        RECT 127.100 3.400 128.900 3.700 ;
        RECT 127.500 3.100 127.800 3.400 ;
        RECT 130.200 3.100 130.600 3.500 ;
        RECT 125.100 1.100 125.700 3.100 ;
        RECT 127.400 1.100 127.800 3.100 ;
        RECT 129.600 2.800 130.600 3.100 ;
        RECT 129.600 1.100 130.000 2.800 ;
        RECT 131.800 1.100 132.200 5.300 ;
        RECT 132.600 1.100 133.000 9.900 ;
        RECT 133.400 8.100 133.800 8.600 ;
        RECT 134.200 8.100 134.600 9.900 ;
        RECT 136.300 9.200 136.900 9.900 ;
        RECT 136.300 8.900 137.000 9.200 ;
        RECT 138.600 8.900 139.000 9.900 ;
        RECT 140.800 9.200 141.200 9.900 ;
        RECT 140.800 8.900 141.800 9.200 ;
        RECT 136.600 8.500 137.000 8.900 ;
        RECT 138.700 8.600 139.000 8.900 ;
        RECT 138.700 8.300 140.100 8.600 ;
        RECT 139.700 8.200 140.100 8.300 ;
        RECT 133.400 7.800 134.600 8.100 ;
        RECT 137.400 7.800 137.800 8.200 ;
        RECT 140.600 7.800 141.000 8.600 ;
        RECT 141.400 8.500 141.800 8.900 ;
        RECT 134.200 7.700 134.600 7.800 ;
        RECT 135.700 7.700 136.100 7.800 ;
        RECT 134.200 7.400 136.100 7.700 ;
        RECT 134.200 5.700 134.600 7.400 ;
        RECT 137.400 7.200 137.700 7.800 ;
        RECT 137.400 7.100 138.100 7.200 ;
        RECT 140.600 7.100 140.900 7.800 ;
        RECT 143.000 7.500 143.400 9.900 ;
        RECT 144.600 7.600 145.000 9.900 ;
        RECT 146.200 7.600 146.600 9.900 ;
        RECT 147.800 7.600 148.200 9.900 ;
        RECT 149.400 7.600 149.800 9.900 ;
        RECT 152.600 7.700 153.000 9.900 ;
        RECT 154.700 9.200 155.300 9.900 ;
        RECT 154.700 8.900 155.400 9.200 ;
        RECT 157.000 8.900 157.400 9.900 ;
        RECT 159.200 9.200 159.600 9.900 ;
        RECT 159.200 8.900 160.200 9.200 ;
        RECT 155.000 8.500 155.400 8.900 ;
        RECT 157.100 8.600 157.400 8.900 ;
        RECT 157.100 8.300 158.500 8.600 ;
        RECT 158.100 8.200 158.500 8.300 ;
        RECT 159.000 8.200 159.400 8.600 ;
        RECT 159.800 8.500 160.200 8.900 ;
        RECT 154.100 7.700 154.500 7.800 ;
        RECT 144.600 7.200 145.500 7.600 ;
        RECT 146.200 7.200 147.300 7.600 ;
        RECT 147.800 7.200 148.900 7.600 ;
        RECT 149.400 7.200 150.600 7.600 ;
        RECT 142.200 7.100 143.000 7.200 ;
        RECT 137.400 6.800 143.000 7.100 ;
        RECT 145.100 6.900 145.500 7.200 ;
        RECT 146.900 6.900 147.300 7.200 ;
        RECT 148.500 6.900 148.900 7.200 ;
        RECT 136.600 6.400 137.000 6.500 ;
        RECT 135.100 6.100 137.000 6.400 ;
        RECT 135.100 6.000 135.500 6.100 ;
        RECT 135.900 5.700 136.300 5.800 ;
        RECT 134.200 5.400 136.300 5.700 ;
        RECT 134.200 1.100 134.600 5.400 ;
        RECT 137.500 5.200 137.800 6.800 ;
        RECT 141.100 6.700 141.500 6.800 ;
        RECT 145.100 6.500 146.400 6.900 ;
        RECT 146.900 6.500 148.100 6.900 ;
        RECT 148.500 6.500 149.800 6.900 ;
        RECT 141.900 6.200 142.300 6.300 ;
        RECT 139.000 6.100 139.400 6.200 ;
        RECT 139.800 6.100 142.300 6.200 ;
        RECT 139.000 5.900 142.300 6.100 ;
        RECT 139.000 5.800 140.200 5.900 ;
        RECT 145.100 5.800 145.500 6.500 ;
        RECT 146.900 5.800 147.300 6.500 ;
        RECT 148.500 5.800 148.900 6.500 ;
        RECT 150.200 5.800 150.600 7.200 ;
        RECT 140.600 5.500 143.400 5.600 ;
        RECT 140.500 5.400 143.400 5.500 ;
        RECT 136.600 4.900 137.800 5.200 ;
        RECT 138.500 5.300 143.400 5.400 ;
        RECT 138.500 5.100 140.900 5.300 ;
        RECT 136.600 4.400 136.900 4.900 ;
        RECT 136.200 4.000 136.900 4.400 ;
        RECT 137.700 4.500 138.100 4.600 ;
        RECT 138.500 4.500 138.800 5.100 ;
        RECT 137.700 4.200 138.800 4.500 ;
        RECT 139.100 4.500 141.800 4.800 ;
        RECT 139.100 4.400 139.500 4.500 ;
        RECT 141.400 4.400 141.800 4.500 ;
        RECT 138.300 3.700 138.700 3.800 ;
        RECT 139.700 3.700 140.100 3.800 ;
        RECT 136.600 3.100 137.000 3.500 ;
        RECT 138.300 3.400 140.100 3.700 ;
        RECT 138.700 3.100 139.000 3.400 ;
        RECT 141.400 3.100 141.800 3.500 ;
        RECT 136.300 1.100 136.900 3.100 ;
        RECT 138.600 1.100 139.000 3.100 ;
        RECT 140.800 2.800 141.800 3.100 ;
        RECT 140.800 1.100 141.200 2.800 ;
        RECT 143.000 1.100 143.400 5.300 ;
        RECT 144.600 5.400 145.500 5.800 ;
        RECT 146.200 5.400 147.300 5.800 ;
        RECT 147.800 5.400 148.900 5.800 ;
        RECT 149.400 5.400 150.600 5.800 ;
        RECT 152.600 7.400 154.500 7.700 ;
        RECT 152.600 5.700 153.000 7.400 ;
        RECT 156.100 7.100 156.500 7.200 ;
        RECT 159.000 7.100 159.300 8.200 ;
        RECT 161.400 7.500 161.800 9.900 ;
        RECT 162.200 7.800 162.600 8.600 ;
        RECT 160.600 7.100 161.400 7.200 ;
        RECT 155.900 6.800 161.400 7.100 ;
        RECT 155.000 6.400 155.400 6.500 ;
        RECT 153.500 6.100 155.400 6.400 ;
        RECT 153.500 6.000 153.900 6.100 ;
        RECT 154.300 5.700 154.700 5.800 ;
        RECT 152.600 5.400 154.700 5.700 ;
        RECT 144.600 1.100 145.000 5.400 ;
        RECT 146.200 1.100 146.600 5.400 ;
        RECT 147.800 1.100 148.200 5.400 ;
        RECT 149.400 1.100 149.800 5.400 ;
        RECT 152.600 1.100 153.000 5.400 ;
        RECT 155.900 5.200 156.200 6.800 ;
        RECT 159.500 6.700 159.900 6.800 ;
        RECT 159.000 6.200 159.400 6.300 ;
        RECT 160.300 6.200 160.700 6.300 ;
        RECT 158.200 5.900 160.700 6.200 ;
        RECT 158.200 5.800 158.600 5.900 ;
        RECT 159.000 5.500 161.800 5.600 ;
        RECT 158.900 5.400 161.800 5.500 ;
        RECT 155.000 4.900 156.200 5.200 ;
        RECT 156.900 5.300 161.800 5.400 ;
        RECT 156.900 5.100 159.300 5.300 ;
        RECT 155.000 4.400 155.300 4.900 ;
        RECT 154.600 4.000 155.300 4.400 ;
        RECT 156.100 4.500 156.500 4.600 ;
        RECT 156.900 4.500 157.200 5.100 ;
        RECT 156.100 4.200 157.200 4.500 ;
        RECT 157.500 4.500 160.200 4.800 ;
        RECT 157.500 4.400 157.900 4.500 ;
        RECT 159.800 4.400 160.200 4.500 ;
        RECT 156.700 3.700 157.100 3.800 ;
        RECT 158.100 3.700 158.500 3.800 ;
        RECT 155.000 3.100 155.400 3.500 ;
        RECT 156.700 3.400 158.500 3.700 ;
        RECT 157.100 3.100 157.400 3.400 ;
        RECT 159.800 3.100 160.200 3.500 ;
        RECT 154.700 1.100 155.300 3.100 ;
        RECT 157.000 1.100 157.400 3.100 ;
        RECT 159.200 2.800 160.200 3.100 ;
        RECT 159.200 1.100 159.600 2.800 ;
        RECT 161.400 1.100 161.800 5.300 ;
        RECT 163.000 1.100 163.400 9.900 ;
        RECT 163.800 7.700 164.200 9.900 ;
        RECT 165.900 9.200 166.500 9.900 ;
        RECT 165.900 8.900 166.600 9.200 ;
        RECT 168.200 8.900 168.600 9.900 ;
        RECT 170.400 9.200 170.800 9.900 ;
        RECT 170.400 8.900 171.400 9.200 ;
        RECT 166.200 8.500 166.600 8.900 ;
        RECT 168.300 8.600 168.600 8.900 ;
        RECT 168.300 8.300 169.700 8.600 ;
        RECT 169.300 8.200 169.700 8.300 ;
        RECT 170.200 8.200 170.600 8.600 ;
        RECT 171.000 8.500 171.400 8.900 ;
        RECT 165.300 7.700 165.700 7.800 ;
        RECT 163.800 7.400 165.700 7.700 ;
        RECT 163.800 5.700 164.200 7.400 ;
        RECT 167.300 7.100 167.700 7.200 ;
        RECT 170.200 7.100 170.500 8.200 ;
        RECT 172.600 7.500 173.000 9.900 ;
        RECT 173.400 7.700 173.800 9.900 ;
        RECT 175.500 9.200 176.100 9.900 ;
        RECT 175.500 8.900 176.200 9.200 ;
        RECT 177.800 8.900 178.200 9.900 ;
        RECT 180.000 9.200 180.400 9.900 ;
        RECT 180.000 8.900 181.000 9.200 ;
        RECT 175.800 8.500 176.200 8.900 ;
        RECT 177.900 8.600 178.200 8.900 ;
        RECT 177.900 8.300 179.300 8.600 ;
        RECT 178.900 8.200 179.300 8.300 ;
        RECT 179.800 8.200 180.200 8.600 ;
        RECT 180.600 8.500 181.000 8.900 ;
        RECT 174.900 7.700 175.300 7.800 ;
        RECT 173.400 7.400 175.300 7.700 ;
        RECT 171.800 7.100 172.600 7.200 ;
        RECT 167.100 6.800 172.600 7.100 ;
        RECT 166.200 6.400 166.600 6.500 ;
        RECT 164.700 6.100 166.600 6.400 ;
        RECT 164.700 6.000 165.100 6.100 ;
        RECT 165.500 5.700 165.900 5.800 ;
        RECT 163.800 5.400 165.900 5.700 ;
        RECT 163.800 1.100 164.200 5.400 ;
        RECT 167.100 5.200 167.400 6.800 ;
        RECT 170.700 6.700 171.100 6.800 ;
        RECT 171.500 6.200 171.900 6.300 ;
        RECT 167.800 6.100 168.200 6.200 ;
        RECT 169.400 6.100 171.900 6.200 ;
        RECT 167.800 5.900 171.900 6.100 ;
        RECT 167.800 5.800 169.800 5.900 ;
        RECT 173.400 5.700 173.800 7.400 ;
        RECT 176.900 7.100 177.300 7.200 ;
        RECT 179.800 7.100 180.100 8.200 ;
        RECT 182.200 7.500 182.600 9.900 ;
        RECT 183.000 7.700 183.400 9.900 ;
        RECT 185.100 9.200 185.700 9.900 ;
        RECT 185.100 8.900 185.800 9.200 ;
        RECT 187.400 8.900 187.800 9.900 ;
        RECT 189.600 9.200 190.000 9.900 ;
        RECT 189.600 8.900 190.600 9.200 ;
        RECT 185.400 8.500 185.800 8.900 ;
        RECT 187.500 8.600 187.800 8.900 ;
        RECT 187.500 8.300 188.900 8.600 ;
        RECT 188.500 8.200 188.900 8.300 ;
        RECT 189.400 8.200 189.800 8.600 ;
        RECT 190.200 8.500 190.600 8.900 ;
        RECT 184.500 7.700 184.900 7.800 ;
        RECT 183.000 7.400 184.900 7.700 ;
        RECT 181.400 7.100 182.200 7.200 ;
        RECT 176.700 6.800 182.200 7.100 ;
        RECT 175.800 6.400 176.200 6.500 ;
        RECT 174.300 6.100 176.200 6.400 ;
        RECT 176.700 6.200 177.000 6.800 ;
        RECT 180.300 6.700 180.700 6.800 ;
        RECT 179.800 6.200 180.200 6.300 ;
        RECT 181.100 6.200 181.500 6.300 ;
        RECT 174.300 6.000 174.700 6.100 ;
        RECT 176.600 5.800 177.000 6.200 ;
        RECT 179.000 5.900 181.500 6.200 ;
        RECT 179.000 5.800 179.400 5.900 ;
        RECT 175.100 5.700 175.500 5.800 ;
        RECT 170.200 5.500 173.000 5.600 ;
        RECT 170.100 5.400 173.000 5.500 ;
        RECT 166.200 4.900 167.400 5.200 ;
        RECT 168.100 5.300 173.000 5.400 ;
        RECT 168.100 5.100 170.500 5.300 ;
        RECT 166.200 4.400 166.500 4.900 ;
        RECT 165.800 4.000 166.500 4.400 ;
        RECT 167.300 4.500 167.700 4.600 ;
        RECT 168.100 4.500 168.400 5.100 ;
        RECT 167.300 4.200 168.400 4.500 ;
        RECT 168.700 4.500 171.400 4.800 ;
        RECT 168.700 4.400 169.100 4.500 ;
        RECT 171.000 4.400 171.400 4.500 ;
        RECT 167.900 3.700 168.300 3.800 ;
        RECT 169.300 3.700 169.700 3.800 ;
        RECT 166.200 3.100 166.600 3.500 ;
        RECT 167.900 3.400 169.700 3.700 ;
        RECT 168.300 3.100 168.600 3.400 ;
        RECT 171.000 3.100 171.400 3.500 ;
        RECT 165.900 1.100 166.500 3.100 ;
        RECT 168.200 1.100 168.600 3.100 ;
        RECT 170.400 2.800 171.400 3.100 ;
        RECT 170.400 1.100 170.800 2.800 ;
        RECT 172.600 1.100 173.000 5.300 ;
        RECT 173.400 5.400 175.500 5.700 ;
        RECT 173.400 1.100 173.800 5.400 ;
        RECT 176.700 5.200 177.000 5.800 ;
        RECT 183.000 5.700 183.400 7.400 ;
        RECT 186.500 7.100 186.900 7.200 ;
        RECT 188.600 7.100 189.000 7.200 ;
        RECT 189.400 7.100 189.700 8.200 ;
        RECT 191.800 7.500 192.200 9.900 ;
        RECT 192.600 7.500 193.000 9.900 ;
        RECT 194.800 9.200 195.200 9.900 ;
        RECT 194.200 8.900 195.200 9.200 ;
        RECT 197.000 8.900 197.400 9.900 ;
        RECT 199.100 9.200 199.700 9.900 ;
        RECT 199.000 8.900 199.700 9.200 ;
        RECT 194.200 8.500 194.600 8.900 ;
        RECT 197.000 8.600 197.300 8.900 ;
        RECT 195.000 8.200 195.400 8.600 ;
        RECT 195.900 8.300 197.300 8.600 ;
        RECT 199.000 8.500 199.400 8.900 ;
        RECT 195.900 8.200 196.300 8.300 ;
        RECT 191.000 7.100 191.800 7.200 ;
        RECT 193.000 7.100 193.800 7.200 ;
        RECT 195.100 7.100 195.400 8.200 ;
        RECT 199.900 7.700 200.300 7.800 ;
        RECT 201.400 7.700 201.800 9.900 ;
        RECT 199.900 7.400 201.800 7.700 ;
        RECT 197.900 7.100 198.300 7.200 ;
        RECT 186.300 6.800 198.500 7.100 ;
        RECT 200.600 6.800 201.000 7.400 ;
        RECT 185.400 6.400 185.800 6.500 ;
        RECT 183.900 6.100 185.800 6.400 ;
        RECT 186.300 6.200 186.600 6.800 ;
        RECT 189.900 6.700 190.300 6.800 ;
        RECT 194.500 6.700 194.900 6.800 ;
        RECT 190.700 6.200 191.100 6.300 ;
        RECT 183.900 6.000 184.300 6.100 ;
        RECT 186.200 5.800 186.600 6.200 ;
        RECT 187.000 6.100 187.400 6.200 ;
        RECT 188.600 6.100 191.100 6.200 ;
        RECT 187.000 5.900 191.100 6.100 ;
        RECT 193.700 6.200 194.100 6.300 ;
        RECT 193.700 5.900 196.200 6.200 ;
        RECT 187.000 5.800 189.000 5.900 ;
        RECT 195.800 5.800 196.200 5.900 ;
        RECT 184.700 5.700 185.100 5.800 ;
        RECT 179.800 5.500 182.600 5.600 ;
        RECT 179.700 5.400 182.600 5.500 ;
        RECT 175.800 4.900 177.000 5.200 ;
        RECT 177.700 5.300 182.600 5.400 ;
        RECT 177.700 5.100 180.100 5.300 ;
        RECT 175.800 4.400 176.100 4.900 ;
        RECT 175.400 4.000 176.100 4.400 ;
        RECT 176.900 4.500 177.300 4.600 ;
        RECT 177.700 4.500 178.000 5.100 ;
        RECT 176.900 4.200 178.000 4.500 ;
        RECT 178.300 4.500 181.000 4.800 ;
        RECT 178.300 4.400 178.700 4.500 ;
        RECT 180.600 4.400 181.000 4.500 ;
        RECT 177.500 3.700 177.900 3.800 ;
        RECT 178.900 3.700 179.300 3.800 ;
        RECT 175.800 3.100 176.200 3.500 ;
        RECT 177.500 3.400 179.300 3.700 ;
        RECT 177.900 3.100 178.200 3.400 ;
        RECT 180.600 3.100 181.000 3.500 ;
        RECT 175.500 1.100 176.100 3.100 ;
        RECT 177.800 1.100 178.200 3.100 ;
        RECT 180.000 2.800 181.000 3.100 ;
        RECT 180.000 1.100 180.400 2.800 ;
        RECT 182.200 1.100 182.600 5.300 ;
        RECT 183.000 5.400 185.100 5.700 ;
        RECT 183.000 1.100 183.400 5.400 ;
        RECT 186.300 5.200 186.600 5.800 ;
        RECT 189.400 5.500 192.200 5.600 ;
        RECT 189.300 5.400 192.200 5.500 ;
        RECT 185.400 4.900 186.600 5.200 ;
        RECT 187.300 5.300 192.200 5.400 ;
        RECT 187.300 5.100 189.700 5.300 ;
        RECT 185.400 4.400 185.700 4.900 ;
        RECT 185.000 4.000 185.700 4.400 ;
        RECT 186.500 4.500 186.900 4.600 ;
        RECT 187.300 4.500 187.600 5.100 ;
        RECT 186.500 4.200 187.600 4.500 ;
        RECT 187.900 4.500 190.600 4.800 ;
        RECT 187.900 4.400 188.300 4.500 ;
        RECT 190.200 4.400 190.600 4.500 ;
        RECT 187.100 3.700 187.500 3.800 ;
        RECT 188.500 3.700 188.900 3.800 ;
        RECT 185.400 3.100 185.800 3.500 ;
        RECT 187.100 3.400 188.900 3.700 ;
        RECT 187.500 3.100 187.800 3.400 ;
        RECT 190.200 3.100 190.600 3.500 ;
        RECT 185.100 1.100 185.700 3.100 ;
        RECT 187.400 1.100 187.800 3.100 ;
        RECT 189.600 2.800 190.600 3.100 ;
        RECT 189.600 1.100 190.000 2.800 ;
        RECT 191.800 1.100 192.200 5.300 ;
        RECT 192.600 5.500 195.400 5.600 ;
        RECT 192.600 5.400 195.500 5.500 ;
        RECT 192.600 5.300 197.500 5.400 ;
        RECT 192.600 1.100 193.000 5.300 ;
        RECT 195.100 5.100 197.500 5.300 ;
        RECT 194.200 4.500 196.900 4.800 ;
        RECT 194.200 4.400 194.600 4.500 ;
        RECT 196.500 4.400 196.900 4.500 ;
        RECT 197.200 4.500 197.500 5.100 ;
        RECT 198.200 5.200 198.500 6.800 ;
        RECT 199.000 6.400 199.400 6.500 ;
        RECT 199.000 6.100 200.900 6.400 ;
        RECT 200.500 6.000 200.900 6.100 ;
        RECT 199.700 5.700 200.100 5.800 ;
        RECT 201.400 5.700 201.800 7.400 ;
        RECT 199.700 5.400 201.800 5.700 ;
        RECT 198.200 4.900 199.400 5.200 ;
        RECT 197.900 4.500 198.300 4.600 ;
        RECT 197.200 4.200 198.300 4.500 ;
        RECT 199.100 4.400 199.400 4.900 ;
        RECT 199.100 4.000 199.800 4.400 ;
        RECT 195.900 3.700 196.300 3.800 ;
        RECT 197.300 3.700 197.700 3.800 ;
        RECT 194.200 3.100 194.600 3.500 ;
        RECT 195.900 3.400 197.700 3.700 ;
        RECT 197.000 3.100 197.300 3.400 ;
        RECT 199.000 3.100 199.400 3.500 ;
        RECT 194.200 2.800 195.200 3.100 ;
        RECT 194.800 1.100 195.200 2.800 ;
        RECT 197.000 1.100 197.400 3.100 ;
        RECT 199.100 1.100 199.700 3.100 ;
        RECT 201.400 1.100 201.800 5.400 ;
        RECT 203.000 1.100 203.400 9.900 ;
      LAYER via1 ;
        RECT 26.200 177.200 26.600 177.600 ;
        RECT 27.800 177.500 28.200 177.900 ;
        RECT 25.400 176.200 25.800 176.600 ;
        RECT 2.200 174.800 2.600 175.200 ;
        RECT 4.600 174.800 5.000 175.200 ;
        RECT 14.200 174.800 14.600 175.200 ;
        RECT 16.600 174.800 17.000 175.200 ;
        RECT 11.000 171.800 11.400 172.200 ;
        RECT 30.200 173.800 30.600 174.200 ;
        RECT 28.600 172.800 29.000 173.200 ;
        RECT 25.400 172.100 25.800 172.500 ;
        RECT 26.200 172.100 26.600 172.500 ;
        RECT 27.000 172.100 27.400 172.500 ;
        RECT 27.800 172.100 28.200 172.500 ;
        RECT 29.400 172.100 29.800 172.500 ;
        RECT 31.000 172.100 31.400 172.500 ;
        RECT 31.800 172.100 32.200 172.500 ;
        RECT 32.600 172.100 33.000 172.500 ;
        RECT 51.000 177.200 51.400 177.600 ;
        RECT 52.600 177.500 53.000 177.900 ;
        RECT 50.200 176.200 50.600 176.600 ;
        RECT 39.800 174.800 40.200 175.200 ;
        RECT 49.400 174.800 49.800 175.200 ;
        RECT 55.000 173.800 55.400 174.200 ;
        RECT 53.400 172.800 53.800 173.200 ;
        RECT 50.200 172.100 50.600 172.500 ;
        RECT 51.000 172.100 51.400 172.500 ;
        RECT 51.800 172.100 52.200 172.500 ;
        RECT 52.600 172.100 53.000 172.500 ;
        RECT 54.200 172.100 54.600 172.500 ;
        RECT 55.800 172.100 56.200 172.500 ;
        RECT 56.600 172.100 57.000 172.500 ;
        RECT 57.400 172.100 57.800 172.500 ;
        RECT 69.400 176.200 69.800 176.600 ;
        RECT 71.000 175.500 71.400 175.900 ;
        RECT 66.200 173.800 66.600 174.200 ;
        RECT 79.000 176.200 79.400 176.600 ;
        RECT 80.600 175.500 81.000 175.900 ;
        RECT 71.000 173.100 71.400 173.500 ;
        RECT 62.200 171.800 62.600 172.200 ;
        RECT 101.400 177.500 101.800 177.900 ;
        RECT 99.800 176.800 100.200 177.200 ;
        RECT 102.200 176.200 102.600 176.600 ;
        RECT 96.600 174.100 97.000 174.500 ;
        RECT 101.400 174.300 101.800 174.700 ;
        RECT 80.600 173.100 81.000 173.500 ;
        RECT 71.800 171.800 72.200 172.200 ;
        RECT 82.200 171.800 82.600 172.200 ;
        RECT 99.000 173.800 99.400 174.200 ;
        RECT 96.600 172.100 97.000 172.500 ;
        RECT 97.400 172.100 97.800 172.500 ;
        RECT 98.200 172.100 98.600 172.500 ;
        RECT 99.800 172.100 100.200 172.500 ;
        RECT 101.400 172.100 101.800 172.500 ;
        RECT 102.200 172.100 102.600 172.500 ;
        RECT 103.000 172.100 103.400 172.500 ;
        RECT 103.800 172.100 104.200 172.500 ;
        RECT 109.400 172.800 109.800 173.200 ;
        RECT 122.200 172.800 122.600 173.200 ;
        RECT 123.000 171.800 123.400 172.200 ;
        RECT 125.400 172.800 125.800 173.200 ;
        RECT 136.600 177.200 137.000 177.600 ;
        RECT 138.200 177.500 138.600 177.900 ;
        RECT 135.800 176.200 136.200 176.600 ;
        RECT 135.000 174.800 135.400 175.200 ;
        RECT 127.000 171.800 127.400 172.200 ;
        RECT 128.600 171.800 129.000 172.200 ;
        RECT 140.600 173.800 141.000 174.200 ;
        RECT 139.000 172.800 139.400 173.200 ;
        RECT 135.800 172.100 136.200 172.500 ;
        RECT 136.600 172.100 137.000 172.500 ;
        RECT 137.400 172.100 137.800 172.500 ;
        RECT 138.200 172.100 138.600 172.500 ;
        RECT 139.800 172.100 140.200 172.500 ;
        RECT 141.400 172.100 141.800 172.500 ;
        RECT 142.200 172.100 142.600 172.500 ;
        RECT 143.000 172.100 143.400 172.500 ;
        RECT 158.200 177.500 158.600 177.900 ;
        RECT 156.600 176.800 157.000 177.200 ;
        RECT 159.000 176.200 159.400 176.600 ;
        RECT 161.400 174.800 161.800 175.200 ;
        RECT 153.400 174.100 153.800 174.500 ;
        RECT 158.200 174.300 158.600 174.700 ;
        RECT 155.800 173.800 156.200 174.200 ;
        RECT 153.400 172.100 153.800 172.500 ;
        RECT 154.200 172.100 154.600 172.500 ;
        RECT 155.000 172.100 155.400 172.500 ;
        RECT 156.600 172.100 157.000 172.500 ;
        RECT 158.200 172.100 158.600 172.500 ;
        RECT 159.000 172.100 159.400 172.500 ;
        RECT 159.800 172.100 160.200 172.500 ;
        RECT 160.600 172.100 161.000 172.500 ;
        RECT 183.000 177.500 183.400 177.900 ;
        RECT 181.400 176.800 181.800 177.200 ;
        RECT 183.800 176.200 184.200 176.600 ;
        RECT 178.200 174.100 178.600 174.500 ;
        RECT 183.000 174.300 183.400 174.700 ;
        RECT 165.400 171.800 165.800 172.200 ;
        RECT 180.600 173.800 181.000 174.200 ;
        RECT 178.200 172.100 178.600 172.500 ;
        RECT 179.000 172.100 179.400 172.500 ;
        RECT 179.800 172.100 180.200 172.500 ;
        RECT 181.400 172.100 181.800 172.500 ;
        RECT 183.000 172.100 183.400 172.500 ;
        RECT 183.800 172.100 184.200 172.500 ;
        RECT 184.600 172.100 185.000 172.500 ;
        RECT 185.400 172.100 185.800 172.500 ;
        RECT 190.200 171.800 190.600 172.200 ;
        RECT 195.000 176.800 195.400 177.200 ;
        RECT 192.600 172.800 193.000 173.200 ;
        RECT 191.800 171.800 192.200 172.200 ;
        RECT 196.600 172.800 197.000 173.200 ;
        RECT 200.600 172.800 201.000 173.200 ;
        RECT 1.400 168.800 1.800 169.200 ;
        RECT 9.400 167.800 9.800 168.200 ;
        RECT 10.200 167.100 10.600 167.500 ;
        RECT 19.000 168.800 19.400 169.200 ;
        RECT 15.800 165.800 16.200 166.200 ;
        RECT 7.000 163.400 7.400 163.800 ;
        RECT 8.600 163.100 9.000 163.500 ;
        RECT 6.200 162.100 6.600 162.500 ;
        RECT 7.000 162.100 7.400 162.500 ;
        RECT 7.800 162.100 8.200 162.500 ;
        RECT 10.200 163.100 10.600 163.500 ;
        RECT 11.800 163.100 12.200 163.500 ;
        RECT 27.000 167.800 27.400 168.200 ;
        RECT 27.800 167.100 28.200 167.500 ;
        RECT 36.600 168.800 37.000 169.200 ;
        RECT 33.400 165.800 33.800 166.200 ;
        RECT 12.600 162.100 13.000 162.500 ;
        RECT 13.400 162.100 13.800 162.500 ;
        RECT 24.600 163.400 25.000 163.800 ;
        RECT 26.200 163.100 26.600 163.500 ;
        RECT 23.800 162.100 24.200 162.500 ;
        RECT 24.600 162.100 25.000 162.500 ;
        RECT 25.400 162.100 25.800 162.500 ;
        RECT 27.800 163.100 28.200 163.500 ;
        RECT 29.400 163.100 29.800 163.500 ;
        RECT 44.600 167.800 45.000 168.200 ;
        RECT 45.400 167.100 45.800 167.500 ;
        RECT 60.600 168.800 61.000 169.200 ;
        RECT 65.400 168.800 65.800 169.200 ;
        RECT 51.000 165.800 51.400 166.200 ;
        RECT 30.200 162.100 30.600 162.500 ;
        RECT 31.000 162.100 31.400 162.500 ;
        RECT 42.200 163.400 42.600 163.800 ;
        RECT 43.800 163.100 44.200 163.500 ;
        RECT 41.400 162.100 41.800 162.500 ;
        RECT 42.200 162.100 42.600 162.500 ;
        RECT 43.000 162.100 43.400 162.500 ;
        RECT 45.400 163.100 45.800 163.500 ;
        RECT 47.000 163.100 47.400 163.500 ;
        RECT 57.400 165.800 57.800 166.200 ;
        RECT 64.600 166.800 65.000 167.200 ;
        RECT 70.200 166.800 70.600 167.200 ;
        RECT 47.800 162.100 48.200 162.500 ;
        RECT 48.600 162.100 49.000 162.500 ;
        RECT 55.800 161.800 56.200 162.200 ;
        RECT 61.400 164.800 61.800 165.200 ;
        RECT 67.000 165.800 67.400 166.200 ;
        RECT 71.800 165.900 72.200 166.300 ;
        RECT 69.400 165.100 69.800 165.500 ;
        RECT 82.200 166.800 82.600 167.200 ;
        RECT 78.200 161.800 78.600 162.200 ;
        RECT 82.200 164.800 82.600 165.200 ;
        RECT 96.600 168.800 97.000 169.200 ;
        RECT 95.800 167.400 96.200 167.800 ;
        RECT 92.600 166.800 93.000 167.200 ;
        RECT 87.000 166.100 87.400 166.500 ;
        RECT 99.000 166.800 99.400 167.200 ;
        RECT 93.400 165.100 93.800 165.500 ;
        RECT 111.800 165.800 112.200 166.200 ;
        RECT 106.200 164.800 106.600 165.200 ;
        RECT 107.000 164.800 107.400 165.200 ;
        RECT 108.600 164.800 109.000 165.200 ;
        RECT 112.600 164.800 113.000 165.200 ;
        RECT 126.200 168.800 126.600 169.200 ;
        RECT 131.000 167.400 131.400 167.800 ;
        RECT 121.400 165.800 121.800 166.200 ;
        RECT 115.800 161.800 116.200 162.200 ;
        RECT 120.600 164.800 121.000 165.200 ;
        RECT 123.800 165.800 124.200 166.200 ;
        RECT 125.400 165.800 125.800 166.200 ;
        RECT 124.600 164.800 125.000 165.200 ;
        RECT 128.600 165.800 129.000 166.200 ;
        RECT 134.200 166.800 134.600 167.200 ;
        RECT 143.800 167.800 144.200 168.200 ;
        RECT 144.600 167.100 145.000 167.500 ;
        RECT 156.600 168.800 157.000 169.200 ;
        RECT 148.600 165.800 149.000 166.200 ;
        RECT 123.000 161.800 123.400 162.200 ;
        RECT 131.800 163.800 132.200 164.200 ;
        RECT 141.400 163.400 141.800 163.800 ;
        RECT 143.000 163.100 143.400 163.500 ;
        RECT 140.600 162.100 141.000 162.500 ;
        RECT 141.400 162.100 141.800 162.500 ;
        RECT 142.200 162.100 142.600 162.500 ;
        RECT 144.600 163.100 145.000 163.500 ;
        RECT 146.200 163.100 146.600 163.500 ;
        RECT 157.400 167.400 157.800 167.800 ;
        RECT 161.400 167.400 161.800 167.800 ;
        RECT 159.000 166.800 159.400 167.200 ;
        RECT 164.600 166.800 165.000 167.200 ;
        RECT 169.400 166.500 169.800 166.900 ;
        RECT 147.000 162.100 147.400 162.500 ;
        RECT 147.800 162.100 148.200 162.500 ;
        RECT 174.200 166.300 174.600 166.700 ;
        RECT 185.400 168.800 185.800 169.200 ;
        RECT 167.000 165.800 167.400 166.200 ;
        RECT 177.400 165.800 177.800 166.200 ;
        RECT 170.200 164.400 170.600 164.800 ;
        RECT 172.600 163.800 173.000 164.200 ;
        RECT 171.000 163.100 171.400 163.500 ;
        RECT 169.400 162.100 169.800 162.500 ;
        RECT 170.200 162.100 170.600 162.500 ;
        RECT 172.600 163.100 173.000 163.500 ;
        RECT 174.200 163.100 174.600 163.500 ;
        RECT 175.000 162.100 175.400 162.500 ;
        RECT 175.800 162.100 176.200 162.500 ;
        RECT 176.600 162.100 177.000 162.500 ;
        RECT 194.200 168.800 194.600 169.200 ;
        RECT 189.400 166.800 189.800 167.200 ;
        RECT 181.400 161.800 181.800 162.200 ;
        RECT 184.600 164.800 185.000 165.200 ;
        RECT 196.600 166.800 197.000 167.200 ;
        RECT 203.800 167.800 204.200 168.200 ;
        RECT 199.800 165.800 200.200 166.200 ;
        RECT 2.200 154.800 2.600 155.200 ;
        RECT 4.600 154.800 5.000 155.200 ;
        RECT 10.200 154.800 10.600 155.200 ;
        RECT 6.200 153.800 6.600 154.200 ;
        RECT 5.400 153.100 5.800 153.500 ;
        RECT 23.800 157.200 24.200 157.600 ;
        RECT 25.400 157.500 25.800 157.900 ;
        RECT 23.000 156.200 23.400 156.600 ;
        RECT 18.100 154.800 18.500 155.200 ;
        RECT 15.000 152.800 15.400 153.200 ;
        RECT 15.800 151.800 16.200 152.200 ;
        RECT 27.800 153.800 28.200 154.200 ;
        RECT 26.200 152.800 26.600 153.200 ;
        RECT 23.000 152.100 23.400 152.500 ;
        RECT 23.800 152.100 24.200 152.500 ;
        RECT 24.600 152.100 25.000 152.500 ;
        RECT 25.400 152.100 25.800 152.500 ;
        RECT 27.000 152.100 27.400 152.500 ;
        RECT 28.600 152.100 29.000 152.500 ;
        RECT 29.400 152.100 29.800 152.500 ;
        RECT 30.200 152.100 30.600 152.500 ;
        RECT 43.800 154.800 44.200 155.200 ;
        RECT 36.600 151.800 37.000 152.200 ;
        RECT 39.800 152.800 40.200 153.200 ;
        RECT 40.600 153.100 41.000 153.500 ;
        RECT 55.000 153.800 55.400 154.200 ;
        RECT 49.400 151.800 49.800 152.200 ;
        RECT 60.600 153.100 61.000 153.500 ;
        RECT 71.000 154.800 71.400 155.200 ;
        RECT 71.800 154.800 72.200 155.200 ;
        RECT 75.000 153.800 75.400 154.200 ;
        RECT 75.800 153.800 76.200 154.200 ;
        RECT 76.600 153.800 77.000 154.200 ;
        RECT 69.400 151.800 69.800 152.200 ;
        RECT 87.000 157.500 87.400 157.900 ;
        RECT 85.400 156.800 85.800 157.200 ;
        RECT 87.800 156.200 88.200 156.600 ;
        RECT 97.400 156.800 97.800 157.200 ;
        RECT 95.800 155.800 96.200 156.200 ;
        RECT 103.800 158.800 104.200 159.200 ;
        RECT 90.200 154.800 90.600 155.200 ;
        RECT 82.200 154.100 82.600 154.500 ;
        RECT 87.000 154.300 87.400 154.700 ;
        RECT 84.600 153.800 85.000 154.200 ;
        RECT 82.200 152.100 82.600 152.500 ;
        RECT 83.000 152.100 83.400 152.500 ;
        RECT 83.800 152.100 84.200 152.500 ;
        RECT 85.400 152.100 85.800 152.500 ;
        RECT 87.000 152.100 87.400 152.500 ;
        RECT 87.800 152.100 88.200 152.500 ;
        RECT 88.600 152.100 89.000 152.500 ;
        RECT 89.400 152.100 89.800 152.500 ;
        RECT 99.000 154.800 99.400 155.200 ;
        RECT 98.200 153.800 98.600 154.200 ;
        RECT 99.800 151.800 100.200 152.200 ;
        RECT 107.000 153.800 107.400 154.200 ;
        RECT 104.600 152.800 105.000 153.200 ;
        RECT 119.800 153.800 120.200 154.200 ;
        RECT 122.200 153.800 122.600 154.200 ;
        RECT 124.600 155.800 125.000 156.200 ;
        RECT 131.000 157.200 131.400 157.600 ;
        RECT 132.600 157.500 133.000 157.900 ;
        RECT 130.200 156.200 130.600 156.600 ;
        RECT 118.200 151.800 118.600 152.200 ;
        RECT 121.400 151.800 121.800 152.200 ;
        RECT 123.800 151.800 124.200 152.200 ;
        RECT 125.400 151.800 125.800 152.200 ;
        RECT 135.000 153.800 135.400 154.200 ;
        RECT 133.400 152.800 133.800 153.200 ;
        RECT 130.200 152.100 130.600 152.500 ;
        RECT 131.000 152.100 131.400 152.500 ;
        RECT 131.800 152.100 132.200 152.500 ;
        RECT 132.600 152.100 133.000 152.500 ;
        RECT 134.200 152.100 134.600 152.500 ;
        RECT 135.800 152.100 136.200 152.500 ;
        RECT 136.600 152.100 137.000 152.500 ;
        RECT 137.400 152.100 137.800 152.500 ;
        RECT 148.600 157.200 149.000 157.600 ;
        RECT 150.200 157.500 150.600 157.900 ;
        RECT 147.800 156.200 148.200 156.600 ;
        RECT 147.000 154.800 147.400 155.200 ;
        RECT 143.000 151.800 143.400 152.200 ;
        RECT 152.600 153.800 153.000 154.200 ;
        RECT 151.000 152.800 151.400 153.200 ;
        RECT 147.800 152.100 148.200 152.500 ;
        RECT 148.600 152.100 149.000 152.500 ;
        RECT 149.400 152.100 149.800 152.500 ;
        RECT 150.200 152.100 150.600 152.500 ;
        RECT 151.800 152.100 152.200 152.500 ;
        RECT 153.400 152.100 153.800 152.500 ;
        RECT 154.200 152.100 154.600 152.500 ;
        RECT 155.000 152.100 155.400 152.500 ;
        RECT 170.200 157.500 170.600 157.900 ;
        RECT 168.600 156.800 169.000 157.200 ;
        RECT 171.000 156.200 171.400 156.600 ;
        RECT 179.800 158.800 180.200 159.200 ;
        RECT 165.400 154.100 165.800 154.500 ;
        RECT 170.200 154.300 170.600 154.700 ;
        RECT 167.800 153.800 168.200 154.200 ;
        RECT 165.400 152.100 165.800 152.500 ;
        RECT 166.200 152.100 166.600 152.500 ;
        RECT 167.000 152.100 167.400 152.500 ;
        RECT 168.600 152.100 169.000 152.500 ;
        RECT 170.200 152.100 170.600 152.500 ;
        RECT 171.000 152.100 171.400 152.500 ;
        RECT 171.800 152.100 172.200 152.500 ;
        RECT 172.600 152.100 173.000 152.500 ;
        RECT 184.600 154.800 185.000 155.200 ;
        RECT 177.400 151.800 177.800 152.200 ;
        RECT 180.600 152.800 181.000 153.200 ;
        RECT 183.000 152.800 183.400 153.200 ;
        RECT 182.200 151.800 182.600 152.200 ;
        RECT 189.400 154.800 189.800 155.200 ;
        RECT 190.200 154.800 190.600 155.200 ;
        RECT 198.200 154.800 198.600 155.200 ;
        RECT 195.800 153.800 196.200 154.200 ;
        RECT 195.000 153.100 195.400 153.500 ;
        RECT 187.800 151.800 188.200 152.200 ;
        RECT 203.800 151.800 204.200 152.200 ;
        RECT 9.400 148.800 9.800 149.200 ;
        RECT 15.000 148.800 15.400 149.200 ;
        RECT 3.000 146.800 3.400 147.200 ;
        RECT 0.600 145.100 1.000 145.500 ;
        RECT 11.800 146.800 12.200 147.200 ;
        RECT 18.200 146.800 18.600 147.200 ;
        RECT 19.800 146.800 20.200 147.200 ;
        RECT 23.000 146.800 23.400 147.200 ;
        RECT 12.600 144.800 13.000 145.200 ;
        RECT 18.200 144.800 18.600 145.200 ;
        RECT 24.600 145.900 25.000 146.300 ;
        RECT 22.200 145.100 22.600 145.500 ;
        RECT 35.800 146.800 36.200 147.200 ;
        RECT 36.600 145.800 37.000 146.200 ;
        RECT 31.000 141.800 31.400 142.200 ;
        RECT 31.800 145.100 32.200 145.500 ;
        RECT 44.600 146.800 45.000 147.200 ;
        RECT 46.200 145.800 46.600 146.200 ;
        RECT 41.400 145.100 41.800 145.500 ;
        RECT 51.800 141.800 52.200 142.200 ;
        RECT 52.600 141.800 53.000 142.200 ;
        RECT 61.400 148.800 61.800 149.200 ;
        RECT 55.800 144.800 56.200 145.200 ;
        RECT 67.000 147.800 67.400 148.200 ;
        RECT 64.600 145.800 65.000 146.200 ;
        RECT 75.800 147.800 76.200 148.200 ;
        RECT 76.600 147.100 77.000 147.500 ;
        RECT 71.800 145.800 72.200 146.200 ;
        RECT 81.400 145.800 81.800 146.200 ;
        RECT 63.800 141.800 64.200 142.200 ;
        RECT 67.800 141.800 68.200 142.200 ;
        RECT 73.400 143.400 73.800 143.800 ;
        RECT 75.000 143.100 75.400 143.500 ;
        RECT 72.600 142.100 73.000 142.500 ;
        RECT 73.400 142.100 73.800 142.500 ;
        RECT 74.200 142.100 74.600 142.500 ;
        RECT 76.600 143.100 77.000 143.500 ;
        RECT 78.200 143.100 78.600 143.500 ;
        RECT 79.000 142.100 79.400 142.500 ;
        RECT 79.800 142.100 80.200 142.500 ;
        RECT 88.600 146.800 89.000 147.200 ;
        RECT 85.400 141.800 85.800 142.200 ;
        RECT 89.400 144.800 89.800 145.200 ;
        RECT 101.400 146.800 101.800 147.200 ;
        RECT 94.200 146.100 94.600 146.500 ;
        RECT 100.600 145.100 101.000 145.500 ;
        RECT 104.600 145.800 105.000 146.200 ;
        RECT 105.400 145.800 105.800 146.200 ;
        RECT 91.800 141.800 92.200 142.200 ;
        RECT 106.200 144.800 106.600 145.200 ;
        RECT 109.400 145.800 109.800 146.200 ;
        RECT 111.800 144.800 112.200 145.200 ;
        RECT 133.400 148.800 133.800 149.200 ;
        RECT 127.000 145.800 127.400 146.200 ;
        RECT 131.800 145.800 132.200 146.200 ;
        RECT 140.600 148.800 141.000 149.200 ;
        RECT 135.000 145.800 135.400 146.200 ;
        RECT 141.400 147.400 141.800 147.800 ;
        RECT 155.000 148.800 155.400 149.200 ;
        RECT 137.400 145.800 137.800 146.200 ;
        RECT 116.600 141.800 117.000 142.200 ;
        RECT 118.200 141.800 118.600 142.200 ;
        RECT 123.000 141.800 123.400 142.200 ;
        RECT 126.200 141.800 126.600 142.200 ;
        RECT 127.800 141.800 128.200 142.200 ;
        RECT 145.400 144.800 145.800 145.200 ;
        RECT 149.400 146.800 149.800 147.200 ;
        RECT 144.600 141.800 145.000 142.200 ;
        RECT 148.600 145.800 149.000 146.200 ;
        RECT 155.800 146.800 156.200 147.200 ;
        RECT 169.400 148.800 169.800 149.200 ;
        RECT 171.000 146.800 171.400 147.200 ;
        RECT 163.800 144.800 164.200 145.200 ;
        RECT 171.000 145.800 171.400 146.200 ;
        RECT 167.000 144.800 167.400 145.200 ;
        RECT 177.400 146.800 177.800 147.200 ;
        RECT 173.400 144.800 173.800 145.200 ;
        RECT 176.600 145.800 177.000 146.200 ;
        RECT 172.600 141.800 173.000 142.200 ;
        RECT 183.800 148.800 184.200 149.200 ;
        RECT 182.200 146.800 182.600 147.200 ;
        RECT 183.000 146.800 183.400 147.200 ;
        RECT 179.800 145.800 180.200 146.200 ;
        RECT 179.000 144.800 179.400 145.200 ;
        RECT 185.400 145.800 185.800 146.200 ;
        RECT 186.200 145.800 186.600 146.200 ;
        RECT 195.800 147.800 196.200 148.200 ;
        RECT 178.200 141.800 178.600 142.200 ;
        RECT 180.600 143.800 181.000 144.200 ;
        RECT 192.600 145.800 193.000 146.200 ;
        RECT 202.200 146.800 202.600 147.200 ;
        RECT 195.000 143.800 195.400 144.200 ;
        RECT 195.800 141.800 196.200 142.200 ;
        RECT 199.800 141.800 200.200 142.200 ;
        RECT 1.400 138.800 1.800 139.200 ;
        RECT 7.000 137.200 7.400 137.600 ;
        RECT 8.600 137.500 9.000 137.900 ;
        RECT 19.000 138.800 19.400 139.200 ;
        RECT 6.200 136.200 6.600 136.600 ;
        RECT 11.000 133.800 11.400 134.200 ;
        RECT 9.400 132.800 9.800 133.200 ;
        RECT 6.200 132.100 6.600 132.500 ;
        RECT 7.000 132.100 7.400 132.500 ;
        RECT 7.800 132.100 8.200 132.500 ;
        RECT 8.600 132.100 9.000 132.500 ;
        RECT 10.200 132.100 10.600 132.500 ;
        RECT 11.800 132.100 12.200 132.500 ;
        RECT 12.600 132.100 13.000 132.500 ;
        RECT 13.400 132.100 13.800 132.500 ;
        RECT 21.400 138.800 21.800 139.200 ;
        RECT 27.000 137.200 27.400 137.600 ;
        RECT 28.600 137.500 29.000 137.900 ;
        RECT 26.200 136.200 26.600 136.600 ;
        RECT 19.800 133.800 20.200 134.200 ;
        RECT 25.400 134.800 25.800 135.200 ;
        RECT 31.000 133.800 31.400 134.200 ;
        RECT 29.400 132.800 29.800 133.200 ;
        RECT 39.000 134.800 39.400 135.200 ;
        RECT 62.200 136.800 62.600 137.200 ;
        RECT 26.200 132.100 26.600 132.500 ;
        RECT 27.000 132.100 27.400 132.500 ;
        RECT 27.800 132.100 28.200 132.500 ;
        RECT 28.600 132.100 29.000 132.500 ;
        RECT 30.200 132.100 30.600 132.500 ;
        RECT 31.800 132.100 32.200 132.500 ;
        RECT 32.600 132.100 33.000 132.500 ;
        RECT 33.400 132.100 33.800 132.500 ;
        RECT 46.200 134.800 46.600 135.200 ;
        RECT 45.400 133.800 45.800 134.200 ;
        RECT 40.600 131.800 41.000 132.200 ;
        RECT 47.000 133.800 47.400 134.200 ;
        RECT 43.000 131.800 43.400 132.200 ;
        RECT 55.800 134.800 56.200 135.200 ;
        RECT 51.800 133.800 52.200 134.200 ;
        RECT 48.600 131.800 49.000 132.200 ;
        RECT 52.600 133.100 53.000 133.500 ;
        RECT 62.200 133.800 62.600 134.200 ;
        RECT 55.000 132.800 55.400 133.200 ;
        RECT 66.200 134.800 66.600 135.200 ;
        RECT 67.000 133.800 67.400 134.200 ;
        RECT 72.600 133.800 73.000 134.200 ;
        RECT 61.400 131.800 61.800 132.200 ;
        RECT 70.200 131.800 70.600 132.200 ;
        RECT 76.600 133.800 77.000 134.200 ;
        RECT 80.600 134.800 81.000 135.200 ;
        RECT 81.400 133.800 81.800 134.200 ;
        RECT 89.400 136.200 89.800 136.600 ;
        RECT 91.000 135.500 91.400 135.900 ;
        RECT 71.800 131.800 72.200 132.200 ;
        RECT 75.000 131.800 75.400 132.200 ;
        RECT 91.800 133.800 92.200 134.200 ;
        RECT 91.000 133.100 91.400 133.500 ;
        RECT 82.200 131.800 82.600 132.200 ;
        RECT 95.800 134.800 96.200 135.200 ;
        RECT 96.600 133.800 97.000 134.200 ;
        RECT 102.200 134.800 102.600 135.200 ;
        RECT 105.400 134.800 105.800 135.200 ;
        RECT 106.200 134.800 106.600 135.200 ;
        RECT 104.600 133.800 105.000 134.200 ;
        RECT 111.000 134.800 111.400 135.200 ;
        RECT 98.200 132.800 98.600 133.200 ;
        RECT 115.000 133.800 115.400 134.200 ;
        RECT 123.000 136.200 123.400 136.600 ;
        RECT 124.600 135.500 125.000 135.900 ;
        RECT 112.600 131.800 113.000 132.200 ;
        RECT 124.600 133.100 125.000 133.500 ;
        RECT 115.800 131.800 116.200 132.200 ;
        RECT 126.200 132.800 126.600 133.200 ;
        RECT 141.400 138.800 141.800 139.200 ;
        RECT 145.400 138.800 145.800 139.200 ;
        RECT 132.600 132.800 133.000 133.200 ;
        RECT 135.000 132.800 135.400 133.200 ;
        RECT 143.000 134.800 143.400 135.200 ;
        RECT 156.600 134.800 157.000 135.200 ;
        RECT 152.600 133.800 153.000 134.200 ;
        RECT 151.800 133.100 152.200 133.500 ;
        RECT 161.400 132.800 161.800 133.200 ;
        RECT 163.000 132.800 163.400 133.200 ;
        RECT 163.800 132.800 164.200 133.200 ;
        RECT 165.400 134.800 165.800 135.200 ;
        RECT 166.200 134.800 166.600 135.200 ;
        RECT 175.800 138.800 176.200 139.200 ;
        RECT 176.600 136.800 177.000 137.200 ;
        RECT 174.200 134.800 174.600 135.200 ;
        RECT 178.200 135.800 178.600 136.200 ;
        RECT 177.400 134.800 177.800 135.200 ;
        RECT 175.000 133.800 175.400 134.200 ;
        RECT 167.800 131.800 168.200 132.200 ;
        RECT 179.000 133.800 179.400 134.200 ;
        RECT 180.600 133.800 181.000 134.200 ;
        RECT 186.200 134.800 186.600 135.200 ;
        RECT 191.000 138.800 191.400 139.200 ;
        RECT 189.400 133.800 189.800 134.200 ;
        RECT 192.600 138.800 193.000 139.200 ;
        RECT 193.400 136.800 193.800 137.200 ;
        RECT 195.000 135.800 195.400 136.200 ;
        RECT 201.400 138.800 201.800 139.200 ;
        RECT 199.800 135.900 200.200 136.300 ;
        RECT 194.200 134.800 194.600 135.200 ;
        RECT 191.800 133.800 192.200 134.200 ;
        RECT 199.800 133.100 200.200 133.500 ;
        RECT 204.600 133.800 205.000 134.200 ;
        RECT 202.200 133.200 202.600 133.600 ;
        RECT 11.000 127.800 11.400 128.200 ;
        RECT 5.400 125.800 5.800 126.200 ;
        RECT 0.600 125.100 1.000 125.500 ;
        RECT 25.400 128.800 25.800 129.200 ;
        RECT 12.600 125.800 13.000 126.200 ;
        RECT 17.400 126.800 17.800 127.200 ;
        RECT 16.600 125.100 17.000 125.500 ;
        RECT 46.200 128.800 46.600 129.200 ;
        RECT 49.400 128.800 49.800 129.200 ;
        RECT 35.800 125.800 36.200 126.200 ;
        RECT 29.400 124.800 29.800 125.200 ;
        RECT 31.800 125.100 32.200 125.500 ;
        RECT 41.400 123.800 41.800 124.200 ;
        RECT 50.200 126.800 50.600 127.200 ;
        RECT 43.000 124.800 43.400 125.200 ;
        RECT 46.200 124.800 46.600 125.200 ;
        RECT 53.400 126.800 53.800 127.200 ;
        RECT 57.400 124.800 57.800 125.200 ;
        RECT 59.000 124.800 59.400 125.200 ;
        RECT 55.000 122.800 55.400 123.200 ;
        RECT 72.600 128.800 73.000 129.200 ;
        RECT 67.800 126.800 68.200 127.200 ;
        RECT 71.000 125.800 71.400 126.200 ;
        RECT 62.200 121.800 62.600 122.200 ;
        RECT 68.600 124.800 69.000 125.200 ;
        RECT 78.200 126.800 78.600 127.200 ;
        RECT 89.400 128.800 89.800 129.200 ;
        RECT 87.800 127.800 88.200 128.200 ;
        RECT 75.000 126.100 75.400 126.500 ;
        RECT 71.800 124.800 72.200 125.200 ;
        RECT 81.400 125.100 81.800 125.500 ;
        RECT 72.600 121.800 73.000 122.200 ;
        RECT 85.400 125.800 85.800 126.200 ;
        RECT 83.800 121.800 84.200 122.200 ;
        RECT 86.200 121.800 86.600 122.200 ;
        RECT 91.800 126.100 92.200 126.500 ;
        RECT 107.000 126.800 107.400 127.200 ;
        RECT 109.400 126.800 109.800 127.200 ;
        RECT 98.200 125.100 98.600 125.500 ;
        RECT 100.600 124.800 101.000 125.200 ;
        RECT 113.400 125.800 113.800 126.200 ;
        RECT 118.200 128.800 118.600 129.200 ;
        RECT 117.400 125.800 117.800 126.200 ;
        RECT 123.800 126.800 124.200 127.200 ;
        RECT 136.600 128.800 137.000 129.200 ;
        RECT 120.600 126.100 121.000 126.500 ;
        RECT 127.000 125.100 127.400 125.500 ;
        RECT 127.800 125.100 128.200 125.500 ;
        RECT 139.000 126.800 139.400 127.200 ;
        RECT 135.000 123.800 135.400 124.200 ;
        RECT 140.600 124.800 141.000 125.200 ;
        RECT 143.800 121.800 144.200 122.200 ;
        RECT 144.600 128.800 145.000 129.200 ;
        RECT 147.000 126.100 147.400 126.500 ;
        RECT 151.000 125.900 151.400 126.300 ;
        RECT 153.400 125.100 153.800 125.500 ;
        RECT 157.400 125.800 157.800 126.200 ;
        RECT 159.800 126.800 160.200 127.200 ;
        RECT 169.400 128.800 169.800 129.200 ;
        RECT 160.600 125.800 161.000 126.200 ;
        RECT 163.000 126.800 163.400 127.200 ;
        RECT 163.800 125.800 164.200 126.200 ;
        RECT 144.600 121.800 145.000 122.200 ;
        RECT 168.600 126.800 169.000 127.200 ;
        RECT 177.400 124.800 177.800 125.200 ;
        RECT 175.800 121.800 176.200 122.200 ;
        RECT 179.800 124.800 180.200 125.200 ;
        RECT 180.600 121.800 181.000 122.200 ;
        RECT 187.000 126.800 187.400 127.200 ;
        RECT 188.600 121.800 189.000 122.200 ;
        RECT 199.000 128.800 199.400 129.200 ;
        RECT 197.400 126.800 197.800 127.200 ;
        RECT 198.200 126.800 198.600 127.200 ;
        RECT 191.000 121.800 191.400 122.200 ;
        RECT 200.600 125.800 201.000 126.200 ;
        RECT 204.600 125.800 205.000 126.200 ;
        RECT 5.400 114.800 5.800 115.200 ;
        RECT 17.400 116.800 17.800 117.200 ;
        RECT 0.600 113.100 1.000 113.500 ;
        RECT 14.200 114.800 14.600 115.200 ;
        RECT 11.000 113.800 11.400 114.200 ;
        RECT 9.400 111.800 9.800 112.200 ;
        RECT 10.200 113.100 10.600 113.500 ;
        RECT 21.400 114.800 21.800 115.200 ;
        RECT 22.200 114.800 22.600 115.200 ;
        RECT 35.800 116.800 36.200 117.200 ;
        RECT 29.400 114.800 29.800 115.200 ;
        RECT 27.000 113.800 27.400 114.200 ;
        RECT 23.800 112.800 24.200 113.200 ;
        RECT 26.200 113.100 26.600 113.500 ;
        RECT 35.800 113.800 36.200 114.200 ;
        RECT 39.800 114.800 40.200 115.200 ;
        RECT 42.200 114.800 42.600 115.200 ;
        RECT 40.600 113.800 41.000 114.200 ;
        RECT 35.000 111.800 35.400 112.200 ;
        RECT 51.000 114.800 51.400 115.200 ;
        RECT 52.600 114.800 53.000 115.200 ;
        RECT 53.400 114.800 53.800 115.200 ;
        RECT 64.600 117.800 65.000 118.200 ;
        RECT 45.400 111.800 45.800 112.200 ;
        RECT 58.200 113.800 58.600 114.200 ;
        RECT 55.000 111.800 55.400 112.200 ;
        RECT 61.400 114.800 61.800 115.200 ;
        RECT 62.200 114.800 62.600 115.200 ;
        RECT 63.000 113.800 63.400 114.200 ;
        RECT 71.800 116.200 72.200 116.600 ;
        RECT 75.000 118.800 75.400 119.200 ;
        RECT 73.400 115.500 73.800 115.900 ;
        RECT 79.000 118.800 79.400 119.200 ;
        RECT 59.000 111.800 59.400 112.200 ;
        RECT 73.400 113.100 73.800 113.500 ;
        RECT 77.400 114.800 77.800 115.200 ;
        RECT 87.000 114.800 87.400 115.200 ;
        RECT 87.800 114.800 88.200 115.200 ;
        RECT 88.600 113.800 89.000 114.200 ;
        RECT 90.200 113.800 90.600 114.200 ;
        RECT 79.000 111.800 79.400 112.200 ;
        RECT 96.600 114.800 97.000 115.200 ;
        RECT 93.400 113.800 93.800 114.200 ;
        RECT 92.600 113.100 93.000 113.500 ;
        RECT 82.200 111.800 82.600 112.200 ;
        RECT 113.400 115.900 113.800 116.300 ;
        RECT 123.000 118.800 123.400 119.200 ;
        RECT 107.800 114.800 108.200 115.200 ;
        RECT 108.600 113.800 109.000 114.200 ;
        RECT 119.000 115.800 119.400 116.200 ;
        RECT 111.800 113.800 112.200 114.200 ;
        RECT 102.200 111.800 102.600 112.200 ;
        RECT 113.400 113.100 113.800 113.500 ;
        RECT 129.400 117.800 129.800 118.200 ;
        RECT 117.400 113.800 117.800 114.200 ;
        RECT 115.800 113.200 116.200 113.600 ;
        RECT 120.600 114.800 121.000 115.200 ;
        RECT 123.800 114.800 124.200 115.200 ;
        RECT 123.800 113.800 124.200 114.200 ;
        RECT 129.400 114.800 129.800 115.200 ;
        RECT 130.200 113.800 130.600 114.200 ;
        RECT 131.000 113.800 131.400 114.200 ;
        RECT 139.800 117.200 140.200 117.600 ;
        RECT 141.400 117.500 141.800 117.900 ;
        RECT 139.000 116.200 139.400 116.600 ;
        RECT 132.600 113.800 133.000 114.200 ;
        RECT 138.200 114.800 138.600 115.200 ;
        RECT 134.200 111.800 134.600 112.200 ;
        RECT 163.000 118.800 163.400 119.200 ;
        RECT 162.200 116.800 162.600 117.200 ;
        RECT 143.800 113.800 144.200 114.200 ;
        RECT 142.200 112.800 142.600 113.200 ;
        RECT 139.000 112.100 139.400 112.500 ;
        RECT 139.800 112.100 140.200 112.500 ;
        RECT 140.600 112.100 141.000 112.500 ;
        RECT 141.400 112.100 141.800 112.500 ;
        RECT 143.000 112.100 143.400 112.500 ;
        RECT 144.600 112.100 145.000 112.500 ;
        RECT 145.400 112.100 145.800 112.500 ;
        RECT 146.200 112.100 146.600 112.500 ;
        RECT 152.600 112.800 153.000 113.200 ;
        RECT 163.800 115.800 164.200 116.200 ;
        RECT 163.000 114.800 163.400 115.200 ;
        RECT 165.400 114.800 165.800 115.200 ;
        RECT 176.600 117.500 177.000 117.900 ;
        RECT 175.000 116.800 175.400 117.200 ;
        RECT 183.800 117.800 184.200 118.200 ;
        RECT 177.400 116.200 177.800 116.600 ;
        RECT 159.000 112.800 159.400 113.200 ;
        RECT 155.800 111.800 156.200 112.200 ;
        RECT 171.800 114.100 172.200 114.500 ;
        RECT 176.600 114.300 177.000 114.700 ;
        RECT 174.200 113.800 174.600 114.200 ;
        RECT 171.800 112.100 172.200 112.500 ;
        RECT 172.600 112.100 173.000 112.500 ;
        RECT 173.400 112.100 173.800 112.500 ;
        RECT 175.000 112.100 175.400 112.500 ;
        RECT 176.600 112.100 177.000 112.500 ;
        RECT 177.400 112.100 177.800 112.500 ;
        RECT 178.200 112.100 178.600 112.500 ;
        RECT 179.000 112.100 179.400 112.500 ;
        RECT 192.600 116.200 193.000 116.600 ;
        RECT 194.200 115.500 194.600 115.900 ;
        RECT 203.800 118.800 204.200 119.200 ;
        RECT 194.200 113.100 194.600 113.500 ;
        RECT 185.400 111.800 185.800 112.200 ;
        RECT 195.000 113.100 195.400 113.500 ;
        RECT 0.600 108.800 1.000 109.200 ;
        RECT 6.200 106.800 6.600 107.200 ;
        RECT 3.000 106.100 3.400 106.500 ;
        RECT 7.000 105.900 7.400 106.300 ;
        RECT 9.400 105.100 9.800 105.500 ;
        RECT 17.400 106.800 17.800 107.200 ;
        RECT 17.400 105.800 17.800 106.200 ;
        RECT 15.000 104.800 15.400 105.200 ;
        RECT 11.000 102.800 11.400 103.200 ;
        RECT 27.800 108.800 28.200 109.200 ;
        RECT 26.200 105.800 26.600 106.200 ;
        RECT 26.200 104.800 26.600 105.200 ;
        RECT 29.400 106.800 29.800 107.200 ;
        RECT 38.200 105.800 38.600 106.200 ;
        RECT 44.600 108.800 45.000 109.200 ;
        RECT 41.400 106.800 41.800 107.200 ;
        RECT 43.800 106.800 44.200 107.200 ;
        RECT 42.200 105.800 42.600 106.200 ;
        RECT 52.600 108.800 53.000 109.200 ;
        RECT 55.000 108.800 55.400 109.200 ;
        RECT 51.000 105.800 51.400 106.200 ;
        RECT 35.800 101.800 36.200 102.200 ;
        RECT 58.200 108.800 58.600 109.200 ;
        RECT 57.400 106.800 57.800 107.200 ;
        RECT 56.600 105.800 57.000 106.200 ;
        RECT 63.800 105.800 64.200 106.200 ;
        RECT 67.000 108.800 67.400 109.200 ;
        RECT 71.800 108.800 72.200 109.200 ;
        RECT 67.800 106.800 68.200 107.200 ;
        RECT 84.600 108.800 85.000 109.200 ;
        RECT 72.600 106.800 73.000 107.200 ;
        RECT 68.600 105.800 69.000 106.200 ;
        RECT 75.000 105.800 75.400 106.200 ;
        RECT 79.800 105.800 80.200 106.200 ;
        RECT 75.800 105.100 76.200 105.500 ;
        RECT 65.400 101.800 65.800 102.200 ;
        RECT 94.200 107.800 94.600 108.200 ;
        RECT 85.400 104.800 85.800 105.200 ;
        RECT 87.800 105.800 88.200 106.200 ;
        RECT 95.800 105.800 96.200 106.200 ;
        RECT 88.600 101.800 89.000 102.200 ;
        RECT 94.200 101.800 94.600 102.200 ;
        RECT 96.600 101.800 97.000 102.200 ;
        RECT 99.800 104.800 100.200 105.200 ;
        RECT 113.400 106.800 113.800 107.200 ;
        RECT 107.800 106.100 108.200 106.500 ;
        RECT 127.000 108.800 127.400 109.200 ;
        RECT 131.000 108.800 131.400 109.200 ;
        RECT 114.200 105.100 114.600 105.500 ;
        RECT 105.400 103.800 105.800 104.200 ;
        RECT 118.200 105.100 118.600 105.500 ;
        RECT 116.600 102.800 117.000 103.200 ;
        RECT 129.400 105.800 129.800 106.200 ;
        RECT 131.800 106.800 132.200 107.200 ;
        RECT 138.200 107.800 138.600 108.200 ;
        RECT 132.600 105.800 133.000 106.200 ;
        RECT 137.400 106.800 137.800 107.200 ;
        RECT 136.600 105.800 137.000 106.200 ;
        RECT 147.800 106.800 148.200 107.200 ;
        RECT 159.800 107.800 160.200 108.200 ;
        RECT 142.200 106.100 142.600 106.500 ;
        RECT 155.800 105.800 156.200 106.200 ;
        RECT 148.600 105.100 149.000 105.500 ;
        RECT 151.000 105.100 151.400 105.500 ;
        RECT 162.200 108.800 162.600 109.200 ;
        RECT 161.400 106.800 161.800 107.200 ;
        RECT 163.800 105.800 164.200 106.200 ;
        RECT 172.600 108.800 173.000 109.200 ;
        RECT 175.800 107.800 176.200 108.200 ;
        RECT 185.400 106.800 185.800 107.200 ;
        RECT 199.000 108.800 199.400 109.200 ;
        RECT 179.800 106.100 180.200 106.500 ;
        RECT 183.800 105.900 184.200 106.300 ;
        RECT 186.200 105.100 186.600 105.500 ;
        RECT 190.200 105.800 190.600 106.200 ;
        RECT 195.800 105.800 196.200 106.200 ;
        RECT 194.200 104.800 194.600 105.200 ;
        RECT 199.800 104.800 200.200 105.200 ;
        RECT 189.400 101.800 189.800 102.200 ;
        RECT 202.200 104.800 202.600 105.200 ;
        RECT 203.000 101.800 203.400 102.200 ;
        RECT 6.200 98.800 6.600 99.200 ;
        RECT 11.800 94.800 12.200 95.200 ;
        RECT 8.600 93.800 9.000 94.200 ;
        RECT 25.400 98.800 25.800 99.200 ;
        RECT 27.000 98.800 27.400 99.200 ;
        RECT 18.200 94.800 18.600 95.200 ;
        RECT 19.000 94.800 19.400 95.200 ;
        RECT 6.200 91.800 6.600 92.200 ;
        RECT 7.800 93.100 8.200 93.500 ;
        RECT 16.600 93.800 17.000 94.200 ;
        RECT 20.600 93.800 21.000 94.200 ;
        RECT 26.200 92.800 26.600 93.200 ;
        RECT 30.200 97.800 30.600 98.200 ;
        RECT 34.200 94.800 34.600 95.200 ;
        RECT 35.000 94.800 35.400 95.200 ;
        RECT 48.600 98.800 49.000 99.200 ;
        RECT 35.800 93.800 36.200 94.200 ;
        RECT 45.400 94.800 45.800 95.200 ;
        RECT 47.800 94.800 48.200 95.200 ;
        RECT 49.400 94.800 49.800 95.200 ;
        RECT 44.600 93.800 45.000 94.200 ;
        RECT 46.200 93.800 46.600 94.200 ;
        RECT 57.400 95.800 57.800 96.200 ;
        RECT 62.200 98.800 62.600 99.200 ;
        RECT 67.000 98.800 67.400 99.200 ;
        RECT 69.400 98.800 69.800 99.200 ;
        RECT 51.000 93.800 51.400 94.200 ;
        RECT 55.800 94.800 56.200 95.200 ;
        RECT 57.400 94.800 57.800 95.200 ;
        RECT 53.400 92.800 53.800 93.200 ;
        RECT 58.200 93.800 58.600 94.200 ;
        RECT 81.400 97.800 81.800 98.200 ;
        RECT 73.400 94.800 73.800 95.200 ;
        RECT 75.000 94.800 75.400 95.200 ;
        RECT 78.200 94.800 78.600 95.200 ;
        RECT 90.200 98.800 90.600 99.200 ;
        RECT 83.000 94.800 83.400 95.200 ;
        RECT 84.600 94.800 85.000 95.200 ;
        RECT 87.000 94.800 87.400 95.200 ;
        RECT 97.400 98.800 97.800 99.200 ;
        RECT 113.400 96.800 113.800 97.200 ;
        RECT 88.600 94.800 89.000 95.200 ;
        RECT 71.800 93.800 72.200 94.200 ;
        RECT 69.400 91.800 69.800 92.200 ;
        RECT 75.800 93.800 76.200 94.200 ;
        RECT 79.000 93.800 79.400 94.200 ;
        RECT 82.200 93.800 82.600 94.200 ;
        RECT 85.400 93.800 85.800 94.200 ;
        RECT 90.200 93.800 90.600 94.200 ;
        RECT 83.000 92.800 83.400 93.200 ;
        RECT 88.600 91.800 89.000 92.200 ;
        RECT 95.800 94.800 96.200 95.200 ;
        RECT 96.600 93.800 97.000 94.200 ;
        RECT 99.000 94.800 99.400 95.200 ;
        RECT 93.400 91.800 93.800 92.200 ;
        RECT 97.400 91.800 97.800 92.200 ;
        RECT 102.200 94.800 102.600 95.200 ;
        RECT 107.800 94.800 108.200 95.200 ;
        RECT 104.600 93.100 105.000 93.500 ;
        RECT 115.000 94.800 115.400 95.200 ;
        RECT 123.800 97.800 124.200 98.200 ;
        RECT 127.800 98.800 128.200 99.200 ;
        RECT 115.800 93.800 116.200 94.200 ;
        RECT 117.400 93.800 117.800 94.200 ;
        RECT 122.200 94.800 122.600 95.200 ;
        RECT 122.200 93.800 122.600 94.200 ;
        RECT 125.400 94.800 125.800 95.200 ;
        RECT 132.600 94.800 133.000 95.200 ;
        RECT 130.200 93.800 130.600 94.200 ;
        RECT 129.400 93.100 129.800 93.500 ;
        RECT 138.200 91.800 138.600 92.200 ;
        RECT 145.400 94.800 145.800 95.200 ;
        RECT 140.600 92.800 141.000 93.200 ;
        RECT 150.200 93.800 150.600 94.200 ;
        RECT 147.000 91.800 147.400 92.200 ;
        RECT 157.400 93.800 157.800 94.200 ;
        RECT 166.200 94.800 166.600 95.200 ;
        RECT 169.400 94.800 169.800 95.200 ;
        RECT 171.800 94.800 172.200 95.200 ;
        RECT 182.200 98.800 182.600 99.200 ;
        RECT 167.000 93.800 167.400 94.200 ;
        RECT 170.200 93.800 170.600 94.200 ;
        RECT 164.600 91.800 165.000 92.200 ;
        RECT 167.800 91.800 168.200 92.200 ;
        RECT 177.400 94.800 177.800 95.200 ;
        RECT 178.200 94.800 178.600 95.200 ;
        RECT 191.000 96.200 191.400 96.600 ;
        RECT 192.600 95.500 193.000 95.900 ;
        RECT 192.600 93.100 193.000 93.500 ;
        RECT 202.200 96.200 202.600 96.600 ;
        RECT 203.800 95.500 204.200 95.900 ;
        RECT 201.400 92.800 201.800 93.200 ;
        RECT 193.400 91.800 193.800 92.200 ;
        RECT 203.800 93.100 204.200 93.500 ;
        RECT 0.600 88.800 1.000 89.200 ;
        RECT 6.200 86.800 6.600 87.200 ;
        RECT 8.600 86.800 9.000 87.200 ;
        RECT 3.000 86.100 3.400 86.500 ;
        RECT 7.000 85.900 7.400 86.300 ;
        RECT 15.800 86.800 16.200 87.200 ;
        RECT 9.400 85.100 9.800 85.500 ;
        RECT 11.800 84.800 12.200 85.200 ;
        RECT 15.800 84.800 16.200 85.200 ;
        RECT 21.400 88.800 21.800 89.200 ;
        RECT 19.000 86.800 19.400 87.200 ;
        RECT 25.400 86.800 25.800 87.200 ;
        RECT 29.400 86.800 29.800 87.200 ;
        RECT 24.600 85.100 25.000 85.500 ;
        RECT 16.600 81.800 17.000 82.200 ;
        RECT 35.800 85.800 36.200 86.200 ;
        RECT 38.200 86.800 38.600 87.200 ;
        RECT 40.600 86.800 41.000 87.200 ;
        RECT 39.000 85.800 39.400 86.200 ;
        RECT 43.800 86.800 44.200 87.200 ;
        RECT 49.400 88.800 49.800 89.200 ;
        RECT 51.800 86.100 52.200 86.500 ;
        RECT 55.800 85.900 56.200 86.300 ;
        RECT 66.200 88.800 66.600 89.200 ;
        RECT 67.800 88.800 68.200 89.200 ;
        RECT 75.000 88.800 75.400 89.200 ;
        RECT 58.200 85.100 58.600 85.500 ;
        RECT 60.600 84.800 61.000 85.200 ;
        RECT 73.400 85.800 73.800 86.200 ;
        RECT 83.800 88.800 84.200 89.200 ;
        RECT 75.800 86.800 76.200 87.200 ;
        RECT 76.600 85.800 77.000 86.200 ;
        RECT 89.400 88.800 89.800 89.200 ;
        RECT 82.200 86.800 82.600 87.200 ;
        RECT 66.200 81.800 66.600 82.200 ;
        RECT 72.600 82.800 73.000 83.200 ;
        RECT 78.200 84.800 78.600 85.200 ;
        RECT 79.800 85.800 80.200 86.200 ;
        RECT 83.000 84.800 83.400 85.200 ;
        RECT 91.800 86.800 92.200 87.200 ;
        RECT 93.400 81.800 93.800 82.200 ;
        RECT 95.800 81.800 96.200 82.200 ;
        RECT 106.200 86.800 106.600 87.200 ;
        RECT 100.600 84.800 101.000 85.200 ;
        RECT 110.200 86.800 110.600 87.200 ;
        RECT 114.200 86.800 114.600 87.200 ;
        RECT 108.600 86.100 109.000 86.500 ;
        RECT 117.400 86.800 117.800 87.200 ;
        RECT 116.600 85.800 117.000 86.200 ;
        RECT 115.000 85.100 115.400 85.500 ;
        RECT 118.200 85.800 118.600 86.200 ;
        RECT 127.000 86.800 127.400 87.200 ;
        RECT 137.400 88.800 137.800 89.200 ;
        RECT 121.400 86.100 121.800 86.500 ;
        RECT 125.400 85.900 125.800 86.300 ;
        RECT 127.800 85.100 128.200 85.500 ;
        RECT 130.200 85.800 130.600 86.200 ;
        RECT 133.400 86.800 133.800 87.200 ;
        RECT 133.400 85.800 133.800 86.200 ;
        RECT 119.000 83.800 119.400 84.200 ;
        RECT 157.400 88.800 157.800 89.200 ;
        RECT 145.400 86.800 145.800 87.200 ;
        RECT 139.800 86.100 140.200 86.500 ;
        RECT 135.800 81.800 136.200 82.200 ;
        RECT 143.800 85.900 144.200 86.300 ;
        RECT 146.200 85.100 146.600 85.500 ;
        RECT 156.600 86.800 157.000 87.200 ;
        RECT 153.400 85.800 153.800 86.200 ;
        RECT 158.200 86.800 158.600 87.200 ;
        RECT 159.000 85.800 159.400 86.200 ;
        RECT 148.600 81.800 149.000 82.200 ;
        RECT 179.800 88.800 180.200 89.200 ;
        RECT 163.800 86.100 164.200 86.500 ;
        RECT 170.200 85.100 170.600 85.500 ;
        RECT 173.400 84.800 173.800 85.200 ;
        RECT 174.200 84.800 174.600 85.200 ;
        RECT 189.400 86.800 189.800 87.200 ;
        RECT 182.200 86.100 182.600 86.500 ;
        RECT 190.200 85.800 190.600 86.200 ;
        RECT 188.600 85.100 189.000 85.500 ;
        RECT 191.000 85.800 191.400 86.200 ;
        RECT 194.200 85.800 194.600 86.200 ;
        RECT 201.400 86.800 201.800 87.200 ;
        RECT 202.200 86.800 202.600 87.200 ;
        RECT 198.200 86.100 198.600 86.500 ;
        RECT 204.600 85.100 205.000 85.500 ;
        RECT 9.400 78.800 9.800 79.200 ;
        RECT 4.600 74.800 5.000 75.200 ;
        RECT 0.600 73.100 1.000 73.500 ;
        RECT 27.800 78.800 28.200 79.200 ;
        RECT 3.000 72.800 3.400 73.200 ;
        RECT 18.200 74.800 18.600 75.200 ;
        RECT 18.200 73.800 18.600 74.200 ;
        RECT 19.000 73.100 19.400 73.500 ;
        RECT 21.400 72.800 21.800 73.200 ;
        RECT 28.600 73.800 29.000 74.200 ;
        RECT 31.000 78.800 31.400 79.200 ;
        RECT 42.200 76.800 42.600 77.200 ;
        RECT 35.800 74.800 36.200 75.200 ;
        RECT 33.400 73.800 33.800 74.200 ;
        RECT 31.800 72.800 32.200 73.200 ;
        RECT 32.600 73.100 33.000 73.500 ;
        RECT 42.200 73.800 42.600 74.200 ;
        RECT 46.200 74.800 46.600 75.200 ;
        RECT 48.600 74.800 49.000 75.200 ;
        RECT 49.400 74.800 49.800 75.200 ;
        RECT 47.000 73.800 47.400 74.200 ;
        RECT 58.200 74.800 58.600 75.200 ;
        RECT 62.200 74.800 62.600 75.200 ;
        RECT 65.400 74.800 65.800 75.200 ;
        RECT 66.200 74.800 66.600 75.200 ;
        RECT 69.400 74.800 69.800 75.200 ;
        RECT 77.400 78.800 77.800 79.200 ;
        RECT 81.400 78.800 81.800 79.200 ;
        RECT 72.600 74.800 73.000 75.200 ;
        RECT 74.200 74.800 74.600 75.200 ;
        RECT 76.600 74.800 77.000 75.200 ;
        RECT 78.200 74.800 78.600 75.200 ;
        RECT 80.600 74.800 81.000 75.200 ;
        RECT 82.200 74.800 82.600 75.200 ;
        RECT 91.800 78.800 92.200 79.200 ;
        RECT 63.000 73.800 63.400 74.200 ;
        RECT 60.600 72.800 61.000 73.200 ;
        RECT 64.600 73.800 65.000 74.200 ;
        RECT 67.800 72.800 68.200 73.200 ;
        RECT 75.000 73.800 75.400 74.200 ;
        RECT 79.000 73.800 79.400 74.200 ;
        RECT 83.000 73.800 83.400 74.200 ;
        RECT 91.000 74.800 91.400 75.200 ;
        RECT 92.600 74.800 93.000 75.200 ;
        RECT 87.800 71.800 88.200 72.200 ;
        RECT 94.200 72.800 94.600 73.200 ;
        RECT 103.800 76.200 104.200 76.600 ;
        RECT 105.400 75.500 105.800 75.900 ;
        RECT 98.200 73.800 98.600 74.200 ;
        RECT 95.800 72.800 96.200 73.200 ;
        RECT 107.800 73.800 108.200 74.200 ;
        RECT 105.400 73.100 105.800 73.500 ;
        RECT 111.800 74.800 112.200 75.200 ;
        RECT 119.000 76.800 119.400 77.200 ;
        RECT 126.200 76.200 126.600 76.600 ;
        RECT 127.800 75.500 128.200 75.900 ;
        RECT 112.600 73.800 113.000 74.200 ;
        RECT 110.200 72.800 110.600 73.200 ;
        RECT 113.400 72.800 113.800 73.200 ;
        RECT 118.200 73.800 118.600 74.200 ;
        RECT 127.800 73.100 128.200 73.500 ;
        RECT 131.000 72.800 131.400 73.200 ;
        RECT 137.400 74.800 137.800 75.200 ;
        RECT 151.000 76.800 151.400 77.200 ;
        RECT 134.200 72.800 134.600 73.200 ;
        RECT 129.400 71.800 129.800 72.200 ;
        RECT 139.000 72.800 139.400 73.200 ;
        RECT 141.400 73.800 141.800 74.200 ;
        RECT 143.000 73.800 143.400 74.200 ;
        RECT 142.200 73.100 142.600 73.500 ;
        RECT 159.800 74.800 160.200 75.200 ;
        RECT 157.400 73.800 157.800 74.200 ;
        RECT 155.000 72.800 155.400 73.200 ;
        RECT 156.600 72.800 157.000 73.200 ;
        RECT 160.600 73.800 161.000 74.200 ;
        RECT 171.000 78.800 171.400 79.200 ;
        RECT 181.400 76.800 181.800 77.200 ;
        RECT 163.000 73.800 163.400 74.200 ;
        RECT 163.800 72.800 164.200 73.200 ;
        RECT 175.800 74.800 176.200 75.200 ;
        RECT 167.000 71.800 167.400 72.200 ;
        RECT 175.800 72.800 176.200 73.200 ;
        RECT 188.600 76.200 189.000 76.600 ;
        RECT 190.200 75.500 190.600 75.900 ;
        RECT 191.000 78.800 191.400 79.200 ;
        RECT 190.200 73.100 190.600 73.500 ;
        RECT 191.800 72.800 192.200 73.200 ;
        RECT 203.000 76.200 203.400 76.600 ;
        RECT 204.600 75.500 205.000 75.900 ;
        RECT 204.600 73.100 205.000 73.500 ;
        RECT 9.400 68.800 9.800 69.200 ;
        RECT 4.600 65.800 5.000 66.200 ;
        RECT 0.600 65.100 1.000 65.500 ;
        RECT 24.600 68.800 25.000 69.200 ;
        RECT 16.600 66.800 17.000 67.200 ;
        RECT 21.400 66.800 21.800 67.200 ;
        RECT 13.400 65.800 13.800 66.200 ;
        RECT 13.400 64.800 13.800 65.200 ;
        RECT 15.800 65.100 16.200 65.500 ;
        RECT 27.000 66.800 27.400 67.200 ;
        RECT 31.800 65.800 32.200 66.200 ;
        RECT 27.800 64.800 28.200 65.200 ;
        RECT 31.000 64.800 31.400 65.200 ;
        RECT 31.800 64.800 32.200 65.200 ;
        RECT 46.200 68.800 46.600 69.200 ;
        RECT 36.600 65.900 37.000 66.300 ;
        RECT 34.200 65.100 34.600 65.500 ;
        RECT 33.400 63.800 33.800 64.200 ;
        RECT 43.000 66.800 43.400 67.200 ;
        RECT 47.800 66.800 48.200 67.200 ;
        RECT 41.400 63.800 41.800 64.200 ;
        RECT 46.200 64.800 46.600 65.200 ;
        RECT 54.200 64.800 54.600 65.200 ;
        RECT 58.200 64.800 58.600 65.200 ;
        RECT 61.400 66.800 61.800 67.200 ;
        RECT 69.400 67.800 69.800 68.200 ;
        RECT 65.400 65.800 65.800 66.200 ;
        RECT 60.600 65.100 61.000 65.500 ;
        RECT 71.800 68.800 72.200 69.200 ;
        RECT 71.000 66.800 71.400 67.200 ;
        RECT 84.600 68.800 85.000 69.200 ;
        RECT 75.000 65.800 75.400 66.200 ;
        RECT 79.000 64.800 79.400 65.200 ;
        RECT 77.400 63.800 77.800 64.200 ;
        RECT 84.600 65.800 85.000 66.200 ;
        RECT 87.800 64.800 88.200 65.200 ;
        RECT 93.400 64.800 93.800 65.200 ;
        RECT 115.800 68.800 116.200 69.200 ;
        RECT 103.000 66.800 103.400 67.200 ;
        RECT 101.400 65.800 101.800 66.200 ;
        RECT 107.000 65.100 107.400 65.500 ;
        RECT 117.400 66.800 117.800 67.200 ;
        RECT 123.000 67.800 123.400 68.200 ;
        RECT 127.800 66.800 128.200 67.200 ;
        RECT 122.200 66.100 122.600 66.500 ;
        RECT 126.200 65.900 126.600 66.300 ;
        RECT 131.000 66.800 131.400 67.200 ;
        RECT 130.200 65.800 130.600 66.200 ;
        RECT 132.600 65.800 133.000 66.200 ;
        RECT 139.800 68.800 140.200 69.200 ;
        RECT 139.000 66.800 139.400 67.200 ;
        RECT 128.600 65.100 129.000 65.500 ;
        RECT 134.200 64.800 134.600 65.200 ;
        RECT 149.400 68.800 149.800 69.200 ;
        RECT 144.600 65.800 145.000 66.200 ;
        RECT 156.600 66.800 157.000 67.200 ;
        RECT 158.200 65.900 158.600 66.300 ;
        RECT 154.200 64.800 154.600 65.200 ;
        RECT 155.800 65.100 156.200 65.500 ;
        RECT 168.600 65.800 169.000 66.200 ;
        RECT 167.800 64.800 168.200 65.200 ;
        RECT 181.400 66.800 181.800 67.200 ;
        RECT 193.400 68.800 193.800 69.200 ;
        RECT 174.200 66.100 174.600 66.500 ;
        RECT 182.200 65.800 182.600 66.200 ;
        RECT 180.600 65.100 181.000 65.500 ;
        RECT 187.000 66.800 187.400 67.200 ;
        RECT 195.000 68.800 195.400 69.200 ;
        RECT 201.400 68.800 201.800 69.200 ;
        RECT 199.800 65.800 200.200 66.200 ;
        RECT 202.200 66.800 202.600 67.200 ;
        RECT 203.000 65.800 203.400 66.200 ;
        RECT 9.400 58.800 9.800 59.200 ;
        RECT 3.800 54.800 4.200 55.200 ;
        RECT 19.000 56.800 19.400 57.200 ;
        RECT 0.600 53.100 1.000 53.500 ;
        RECT 14.200 54.800 14.600 55.200 ;
        RECT 11.000 53.800 11.400 54.200 ;
        RECT 3.000 52.800 3.400 53.200 ;
        RECT 9.400 51.800 9.800 52.200 ;
        RECT 10.200 53.100 10.600 53.500 ;
        RECT 35.000 56.800 35.400 57.200 ;
        RECT 29.400 54.800 29.800 55.200 ;
        RECT 24.600 53.800 25.000 54.200 ;
        RECT 25.400 53.100 25.800 53.500 ;
        RECT 27.800 52.800 28.200 53.200 ;
        RECT 39.000 54.800 39.400 55.200 ;
        RECT 41.400 54.800 41.800 55.200 ;
        RECT 52.600 56.800 53.000 57.200 ;
        RECT 47.000 54.800 47.400 55.200 ;
        RECT 39.800 53.800 40.200 54.200 ;
        RECT 44.600 53.800 45.000 54.200 ;
        RECT 43.800 53.100 44.200 53.500 ;
        RECT 55.800 54.800 56.200 55.200 ;
        RECT 62.200 58.800 62.600 59.200 ;
        RECT 75.800 57.800 76.200 58.200 ;
        RECT 55.000 53.800 55.400 54.200 ;
        RECT 62.200 54.800 62.600 55.200 ;
        RECT 70.200 54.800 70.600 55.200 ;
        RECT 59.800 53.800 60.200 54.200 ;
        RECT 63.000 53.800 63.400 54.200 ;
        RECT 67.000 53.100 67.400 53.500 ;
        RECT 77.400 54.800 77.800 55.200 ;
        RECT 87.000 58.800 87.400 59.200 ;
        RECT 81.400 53.800 81.800 54.200 ;
        RECT 87.000 54.800 87.400 55.200 ;
        RECT 89.400 54.800 89.800 55.200 ;
        RECT 107.000 58.800 107.400 59.200 ;
        RECT 83.000 52.800 83.400 53.200 ;
        RECT 87.800 53.800 88.200 54.200 ;
        RECT 91.800 53.800 92.200 54.200 ;
        RECT 93.400 53.800 93.800 54.200 ;
        RECT 94.200 53.100 94.600 53.500 ;
        RECT 107.800 53.800 108.200 54.200 ;
        RECT 103.000 51.800 103.400 52.200 ;
        RECT 119.000 56.800 119.400 57.200 ;
        RECT 110.200 53.800 110.600 54.200 ;
        RECT 114.200 54.800 114.600 55.200 ;
        RECT 115.000 53.800 115.400 54.200 ;
        RECT 126.200 56.200 126.600 56.600 ;
        RECT 127.800 55.500 128.200 55.900 ;
        RECT 129.400 54.800 129.800 55.200 ;
        RECT 130.200 54.800 130.600 55.200 ;
        RECT 147.000 58.800 147.400 59.200 ;
        RECT 112.600 51.800 113.000 52.200 ;
        RECT 117.400 51.800 117.800 52.200 ;
        RECT 127.800 53.100 128.200 53.500 ;
        RECT 133.400 53.800 133.800 54.200 ;
        RECT 135.000 53.800 135.400 54.200 ;
        RECT 134.200 53.100 134.600 53.500 ;
        RECT 141.400 53.800 141.800 54.200 ;
        RECT 154.200 56.200 154.600 56.600 ;
        RECT 155.800 55.500 156.200 55.900 ;
        RECT 145.400 51.800 145.800 52.200 ;
        RECT 156.600 53.800 157.000 54.200 ;
        RECT 155.800 53.100 156.200 53.500 ;
        RECT 167.000 56.200 167.400 56.600 ;
        RECT 168.600 55.500 169.000 55.900 ;
        RECT 169.400 54.800 169.800 55.200 ;
        RECT 170.200 54.800 170.600 55.200 ;
        RECT 176.600 58.800 177.000 59.200 ;
        RECT 173.400 54.800 173.800 55.200 ;
        RECT 168.600 53.100 169.000 53.500 ;
        RECT 171.800 52.800 172.200 53.200 ;
        RECT 179.000 54.800 179.400 55.200 ;
        RECT 179.800 53.800 180.200 54.200 ;
        RECT 181.400 53.800 181.800 54.200 ;
        RECT 180.600 53.100 181.000 53.500 ;
        RECT 191.000 58.800 191.400 59.200 ;
        RECT 192.600 58.800 193.000 59.200 ;
        RECT 195.800 51.800 196.200 52.200 ;
        RECT 199.000 52.800 199.400 53.200 ;
        RECT 203.000 51.800 203.400 52.200 ;
        RECT 6.200 48.800 6.600 49.200 ;
        RECT 11.000 48.800 11.400 49.200 ;
        RECT 9.400 45.800 9.800 46.200 ;
        RECT 12.600 46.800 13.000 47.200 ;
        RECT 12.600 45.800 13.000 46.200 ;
        RECT 19.000 46.800 19.400 47.200 ;
        RECT 22.200 46.800 22.600 47.200 ;
        RECT 15.000 44.800 15.400 45.200 ;
        RECT 33.400 48.800 33.800 49.200 ;
        RECT 25.400 46.800 25.800 47.200 ;
        RECT 27.800 46.800 28.200 47.200 ;
        RECT 27.000 45.900 27.400 46.300 ;
        RECT 22.200 44.800 22.600 45.200 ;
        RECT 24.600 45.100 25.000 45.500 ;
        RECT 36.600 46.800 37.000 47.200 ;
        RECT 56.600 48.800 57.000 49.200 ;
        RECT 42.200 45.900 42.600 46.300 ;
        RECT 37.400 44.800 37.800 45.200 ;
        RECT 39.800 45.100 40.200 45.500 ;
        RECT 59.000 48.800 59.400 49.200 ;
        RECT 53.400 44.800 53.800 45.200 ;
        RECT 61.400 46.800 61.800 47.200 ;
        RECT 56.600 44.800 57.000 45.200 ;
        RECT 65.400 45.800 65.800 46.200 ;
        RECT 60.600 45.100 61.000 45.500 ;
        RECT 71.000 46.800 71.400 47.200 ;
        RECT 75.000 45.800 75.400 46.200 ;
        RECT 69.400 41.800 69.800 42.200 ;
        RECT 70.200 45.100 70.600 45.500 ;
        RECT 90.200 48.800 90.600 49.200 ;
        RECT 80.600 45.800 81.000 46.200 ;
        RECT 82.200 45.800 82.600 46.200 ;
        RECT 89.400 46.800 89.800 47.200 ;
        RECT 86.200 45.800 86.600 46.200 ;
        RECT 94.200 48.800 94.600 49.200 ;
        RECT 104.600 48.800 105.000 49.200 ;
        RECT 95.800 46.800 96.200 47.200 ;
        RECT 94.200 44.800 94.600 45.200 ;
        RECT 107.800 48.800 108.200 49.200 ;
        RECT 100.600 46.800 101.000 47.200 ;
        RECT 103.800 46.800 104.200 47.200 ;
        RECT 110.200 48.800 110.600 49.200 ;
        RECT 107.000 46.800 107.400 47.200 ;
        RECT 111.000 46.800 111.400 47.200 ;
        RECT 111.800 45.800 112.200 46.200 ;
        RECT 115.800 45.800 116.200 46.200 ;
        RECT 126.200 46.800 126.600 47.200 ;
        RECT 134.200 48.800 134.600 49.200 ;
        RECT 120.600 46.100 121.000 46.500 ;
        RECT 127.000 45.100 127.400 45.500 ;
        RECT 133.400 45.800 133.800 46.200 ;
        RECT 139.800 46.800 140.200 47.200 ;
        RECT 136.600 46.100 137.000 46.500 ;
        RECT 131.800 41.800 132.200 42.200 ;
        RECT 140.600 45.900 141.000 46.300 ;
        RECT 143.000 45.100 143.400 45.500 ;
        RECT 145.400 45.800 145.800 46.200 ;
        RECT 147.800 46.800 148.200 47.200 ;
        RECT 148.600 45.800 149.000 46.200 ;
        RECT 163.000 48.800 163.400 49.200 ;
        RECT 162.200 46.800 162.600 47.200 ;
        RECT 155.000 41.800 155.400 42.200 ;
        RECT 159.800 45.800 160.200 46.200 ;
        RECT 159.000 41.800 159.400 42.200 ;
        RECT 167.000 45.800 167.400 46.200 ;
        RECT 170.200 44.800 170.600 45.200 ;
        RECT 168.600 41.800 169.000 42.200 ;
        RECT 171.000 41.800 171.400 42.200 ;
        RECT 173.400 41.800 173.800 42.200 ;
        RECT 175.000 45.100 175.400 45.500 ;
        RECT 185.400 45.800 185.800 46.200 ;
        RECT 191.800 46.800 192.200 47.200 ;
        RECT 190.200 45.800 190.600 46.200 ;
        RECT 195.800 45.800 196.200 46.200 ;
        RECT 191.000 45.100 191.400 45.500 ;
        RECT 198.200 43.800 198.600 44.200 ;
        RECT 201.400 48.800 201.800 49.200 ;
        RECT 204.600 45.800 205.000 46.200 ;
        RECT 11.000 38.800 11.400 39.200 ;
        RECT 0.600 32.800 1.000 33.200 ;
        RECT 5.400 34.800 5.800 35.200 ;
        RECT 3.000 33.800 3.400 34.200 ;
        RECT 2.200 33.100 2.600 33.500 ;
        RECT 15.000 34.800 15.400 35.200 ;
        RECT 15.800 34.800 16.200 35.200 ;
        RECT 18.200 34.800 18.600 35.200 ;
        RECT 19.000 34.800 19.400 35.200 ;
        RECT 31.800 36.800 32.200 37.200 ;
        RECT 22.200 34.800 22.600 35.200 ;
        RECT 27.000 34.800 27.400 35.200 ;
        RECT 16.600 32.800 17.000 33.200 ;
        RECT 23.000 33.100 23.400 33.500 ;
        RECT 33.400 34.800 33.800 35.200 ;
        RECT 34.200 34.800 34.600 35.200 ;
        RECT 35.800 33.800 36.200 34.200 ;
        RECT 20.600 31.800 21.000 32.200 ;
        RECT 25.400 32.800 25.800 33.200 ;
        RECT 38.200 32.800 38.600 33.200 ;
        RECT 39.000 31.800 39.400 32.200 ;
        RECT 43.800 34.800 44.200 35.200 ;
        RECT 53.400 38.800 53.800 39.200 ;
        RECT 58.200 38.800 58.600 39.200 ;
        RECT 41.400 31.800 41.800 32.200 ;
        RECT 63.000 35.800 63.400 36.200 ;
        RECT 61.400 34.800 61.800 35.200 ;
        RECT 54.200 32.800 54.600 33.200 ;
        RECT 56.600 32.800 57.000 33.200 ;
        RECT 61.400 33.800 61.800 34.200 ;
        RECT 64.600 34.800 65.000 35.200 ;
        RECT 66.200 34.800 66.600 35.200 ;
        RECT 67.000 34.800 67.400 35.200 ;
        RECT 75.000 38.800 75.400 39.200 ;
        RECT 79.800 38.800 80.200 39.200 ;
        RECT 70.200 33.800 70.600 34.200 ;
        RECT 73.400 34.800 73.800 35.200 ;
        RECT 82.200 34.800 82.600 35.200 ;
        RECT 84.600 34.800 85.000 35.200 ;
        RECT 77.400 33.800 77.800 34.200 ;
        RECT 71.800 31.800 72.200 32.200 ;
        RECT 78.200 32.800 78.600 33.200 ;
        RECT 83.000 33.800 83.400 34.200 ;
        RECT 86.200 33.800 86.600 34.200 ;
        RECT 89.400 38.800 89.800 39.200 ;
        RECT 96.600 36.200 97.000 36.600 ;
        RECT 104.600 38.800 105.000 39.200 ;
        RECT 98.200 35.500 98.600 35.900 ;
        RECT 103.800 34.800 104.200 35.200 ;
        RECT 105.400 34.800 105.800 35.200 ;
        RECT 110.200 34.800 110.600 35.200 ;
        RECT 111.000 34.800 111.400 35.200 ;
        RECT 98.200 33.100 98.600 33.500 ;
        RECT 100.600 32.800 101.000 33.200 ;
        RECT 115.800 33.800 116.200 34.200 ;
        RECT 113.400 31.800 113.800 32.200 ;
        RECT 123.800 36.200 124.200 36.600 ;
        RECT 125.400 35.500 125.800 35.900 ;
        RECT 125.400 33.100 125.800 33.500 ;
        RECT 126.200 32.800 126.600 33.200 ;
        RECT 132.600 34.800 133.000 35.200 ;
        RECT 137.400 36.800 137.800 37.200 ;
        RECT 133.400 34.800 133.800 35.200 ;
        RECT 135.000 34.800 135.400 35.200 ;
        RECT 135.800 34.800 136.200 35.200 ;
        RECT 129.400 31.800 129.800 32.200 ;
        RECT 145.400 36.200 145.800 36.600 ;
        RECT 147.000 35.500 147.400 35.900 ;
        RECT 148.600 38.800 149.000 39.200 ;
        RECT 156.600 38.800 157.000 39.200 ;
        RECT 147.000 33.100 147.400 33.500 ;
        RECT 165.400 36.200 165.800 36.600 ;
        RECT 167.000 35.500 167.400 35.900 ;
        RECT 167.000 33.100 167.400 33.500 ;
        RECT 167.800 32.800 168.200 33.200 ;
        RECT 173.400 34.800 173.800 35.200 ;
        RECT 174.200 34.800 174.600 35.200 ;
        RECT 179.000 35.800 179.400 36.200 ;
        RECT 171.000 31.800 171.400 32.200 ;
        RECT 177.400 33.800 177.800 34.200 ;
        RECT 179.000 32.800 179.400 33.200 ;
        RECT 179.800 32.800 180.200 33.200 ;
        RECT 192.600 36.200 193.000 36.600 ;
        RECT 194.200 35.500 194.600 35.900 ;
        RECT 195.000 38.800 195.400 39.200 ;
        RECT 183.000 31.800 183.400 32.200 ;
        RECT 202.200 36.200 202.600 36.600 ;
        RECT 203.800 35.500 204.200 35.900 ;
        RECT 194.200 33.100 194.600 33.500 ;
        RECT 203.800 33.100 204.200 33.500 ;
        RECT 0.600 28.800 1.000 29.200 ;
        RECT 6.200 26.800 6.600 27.200 ;
        RECT 10.200 28.800 10.600 29.200 ;
        RECT 3.000 26.100 3.400 26.500 ;
        RECT 7.000 25.900 7.400 26.300 ;
        RECT 28.600 28.800 29.000 29.200 ;
        RECT 20.600 26.800 21.000 27.200 ;
        RECT 25.400 26.800 25.800 27.200 ;
        RECT 12.600 26.100 13.000 26.500 ;
        RECT 16.600 25.900 17.000 26.300 ;
        RECT 9.400 25.100 9.800 25.500 ;
        RECT 19.000 25.100 19.400 25.500 ;
        RECT 19.800 25.100 20.200 25.500 ;
        RECT 43.800 28.800 44.200 29.200 ;
        RECT 35.800 26.800 36.200 27.200 ;
        RECT 31.000 24.800 31.400 25.200 ;
        RECT 35.000 25.100 35.400 25.500 ;
        RECT 59.000 28.800 59.400 29.200 ;
        RECT 47.800 24.800 48.200 25.200 ;
        RECT 54.200 25.800 54.600 26.200 ;
        RECT 69.400 28.800 69.800 29.200 ;
        RECT 59.800 26.800 60.200 27.200 ;
        RECT 86.200 28.800 86.600 29.200 ;
        RECT 57.400 24.800 57.800 25.200 ;
        RECT 60.600 25.800 61.000 26.200 ;
        RECT 63.000 25.800 63.400 26.200 ;
        RECT 66.200 25.800 66.600 26.200 ;
        RECT 65.400 24.800 65.800 25.200 ;
        RECT 72.600 25.800 73.000 26.200 ;
        RECT 74.200 25.800 74.600 26.200 ;
        RECT 69.400 24.800 69.800 25.200 ;
        RECT 71.800 24.800 72.200 25.200 ;
        RECT 79.800 24.800 80.200 25.200 ;
        RECT 93.400 26.800 93.800 27.200 ;
        RECT 105.400 28.800 105.800 29.200 ;
        RECT 86.200 24.800 86.600 25.200 ;
        RECT 90.200 25.800 90.600 26.200 ;
        RECT 97.400 25.800 97.800 26.200 ;
        RECT 89.400 21.800 89.800 22.200 ;
        RECT 94.200 24.800 94.600 25.200 ;
        RECT 97.400 24.800 97.800 25.200 ;
        RECT 101.400 25.800 101.800 26.200 ;
        RECT 127.800 28.800 128.200 29.200 ;
        RECT 107.000 25.800 107.400 26.200 ;
        RECT 109.400 25.800 109.800 26.200 ;
        RECT 111.800 26.800 112.200 27.200 ;
        RECT 124.600 26.800 125.000 27.200 ;
        RECT 127.000 26.800 127.400 27.200 ;
        RECT 112.600 25.800 113.000 26.200 ;
        RECT 100.600 21.800 101.000 22.200 ;
        RECT 110.200 21.800 110.600 22.200 ;
        RECT 119.000 25.800 119.400 26.200 ;
        RECT 132.600 26.800 133.000 27.200 ;
        RECT 118.200 21.800 118.600 22.200 ;
        RECT 125.400 24.800 125.800 25.200 ;
        RECT 140.600 26.800 141.000 27.200 ;
        RECT 135.000 26.100 135.400 26.500 ;
        RECT 141.400 25.100 141.800 25.500 ;
        RECT 144.600 28.800 145.000 29.200 ;
        RECT 143.800 25.800 144.200 26.200 ;
        RECT 157.400 28.800 157.800 29.200 ;
        RECT 156.600 26.800 157.000 27.200 ;
        RECT 147.000 26.100 147.400 26.500 ;
        RECT 148.600 25.800 149.000 26.200 ;
        RECT 151.000 25.900 151.400 26.300 ;
        RECT 155.800 25.800 156.200 26.200 ;
        RECT 164.600 28.800 165.000 29.200 ;
        RECT 167.800 28.800 168.200 29.200 ;
        RECT 153.400 25.100 153.800 25.500 ;
        RECT 163.000 26.800 163.400 27.200 ;
        RECT 160.600 25.800 161.000 26.200 ;
        RECT 162.200 25.800 162.600 26.200 ;
        RECT 163.800 25.800 164.200 26.200 ;
        RECT 167.000 25.800 167.400 26.200 ;
        RECT 175.800 26.800 176.200 27.200 ;
        RECT 170.200 26.100 170.600 26.500 ;
        RECT 191.800 28.800 192.200 29.200 ;
        RECT 179.800 26.100 180.200 26.500 ;
        RECT 176.600 25.100 177.000 25.500 ;
        RECT 186.200 25.100 186.600 25.500 ;
        RECT 190.200 25.800 190.600 26.200 ;
        RECT 189.400 21.800 189.800 22.200 ;
        RECT 193.400 27.800 193.800 28.200 ;
        RECT 198.200 25.800 198.600 26.200 ;
        RECT 24.600 16.800 25.000 17.200 ;
        RECT 5.400 14.800 5.800 15.200 ;
        RECT 0.600 13.100 1.000 13.500 ;
        RECT 10.200 13.800 10.600 14.200 ;
        RECT 19.000 14.800 19.400 15.200 ;
        RECT 11.800 12.800 12.200 13.200 ;
        RECT 15.000 12.800 15.400 13.200 ;
        RECT 15.800 13.100 16.200 13.500 ;
        RECT 26.200 14.800 26.600 15.200 ;
        RECT 27.000 14.800 27.400 15.200 ;
        RECT 31.800 14.800 32.200 15.200 ;
        RECT 30.200 13.800 30.600 14.200 ;
        RECT 37.400 18.800 37.800 19.200 ;
        RECT 35.800 13.800 36.200 14.200 ;
        RECT 33.400 11.800 33.800 12.200 ;
        RECT 36.600 12.800 37.000 13.200 ;
        RECT 49.400 17.800 49.800 18.200 ;
        RECT 43.800 14.800 44.200 15.200 ;
        RECT 40.600 13.100 41.000 13.500 ;
        RECT 39.800 11.800 40.200 12.200 ;
        RECT 52.600 14.800 53.000 15.200 ;
        RECT 53.400 14.800 53.800 15.200 ;
        RECT 59.000 18.800 59.400 19.200 ;
        RECT 62.200 18.800 62.600 19.200 ;
        RECT 59.800 14.800 60.200 15.200 ;
        RECT 56.600 13.800 57.000 14.200 ;
        RECT 57.400 12.800 57.800 13.200 ;
        RECT 69.400 16.200 69.800 16.600 ;
        RECT 79.800 18.800 80.200 19.200 ;
        RECT 71.000 15.500 71.400 15.900 ;
        RECT 72.600 14.800 73.000 15.200 ;
        RECT 75.800 14.800 76.200 15.200 ;
        RECT 83.000 18.800 83.400 19.200 ;
        RECT 79.000 14.800 79.400 15.200 ;
        RECT 61.400 12.800 61.800 13.200 ;
        RECT 81.400 14.800 81.800 15.200 ;
        RECT 71.000 13.100 71.400 13.500 ;
        RECT 81.400 13.800 81.800 14.200 ;
        RECT 74.200 11.800 74.600 12.200 ;
        RECT 82.200 12.800 82.600 13.200 ;
        RECT 83.800 13.800 84.200 14.200 ;
        RECT 87.800 14.800 88.200 15.200 ;
        RECT 94.200 14.800 94.600 15.200 ;
        RECT 88.600 13.800 89.000 14.200 ;
        RECT 89.400 13.100 89.800 13.500 ;
        RECT 86.200 11.800 86.600 12.200 ;
        RECT 91.800 12.800 92.200 13.200 ;
        RECT 98.200 12.800 98.600 13.200 ;
        RECT 99.000 18.800 99.400 19.200 ;
        RECT 104.600 18.800 105.000 19.200 ;
        RECT 99.800 12.800 100.200 13.200 ;
        RECT 100.600 12.800 101.000 13.200 ;
        RECT 111.800 16.200 112.200 16.600 ;
        RECT 113.400 15.500 113.800 15.900 ;
        RECT 114.200 13.800 114.600 14.200 ;
        RECT 113.400 13.100 113.800 13.500 ;
        RECT 118.200 14.800 118.600 15.200 ;
        RECT 130.200 18.800 130.600 19.200 ;
        RECT 119.000 13.800 119.400 14.200 ;
        RECT 120.600 13.800 121.000 14.200 ;
        RECT 119.800 13.100 120.200 13.500 ;
        RECT 136.600 14.800 137.000 15.200 ;
        RECT 137.400 14.800 137.800 15.200 ;
        RECT 147.000 17.800 147.400 18.200 ;
        RECT 141.400 14.800 141.800 15.200 ;
        RECT 141.400 12.800 141.800 13.200 ;
        RECT 144.600 12.800 145.000 13.200 ;
        RECT 139.000 11.800 139.400 12.200 ;
        RECT 154.200 16.200 154.600 16.600 ;
        RECT 155.800 15.500 156.200 15.900 ;
        RECT 155.800 13.100 156.200 13.500 ;
        RECT 196.600 18.800 197.000 19.200 ;
        RECT 163.800 12.800 164.200 13.200 ;
        RECT 175.800 14.800 176.200 15.200 ;
        RECT 161.400 11.800 161.800 12.200 ;
        RECT 167.000 11.800 167.400 12.200 ;
        RECT 176.600 12.800 177.000 13.200 ;
        RECT 182.200 12.800 182.600 13.200 ;
        RECT 199.800 18.800 200.200 19.200 ;
        RECT 188.600 13.800 189.000 14.200 ;
        RECT 179.800 11.800 180.200 12.200 ;
        RECT 185.400 11.800 185.800 12.200 ;
        RECT 187.800 13.100 188.200 13.500 ;
        RECT 197.400 14.800 197.800 15.200 ;
        RECT 200.600 12.800 201.000 13.200 ;
        RECT 6.200 8.800 6.600 9.200 ;
        RECT 14.200 6.800 14.600 7.200 ;
        RECT 15.800 6.800 16.200 7.200 ;
        RECT 24.600 7.800 25.000 8.200 ;
        RECT 15.000 5.100 15.400 5.500 ;
        RECT 26.200 5.800 26.600 6.200 ;
        RECT 39.000 8.800 39.400 9.200 ;
        RECT 28.600 6.800 29.000 7.200 ;
        RECT 31.000 6.800 31.400 7.200 ;
        RECT 43.000 8.800 43.400 9.200 ;
        RECT 29.400 5.800 29.800 6.200 ;
        RECT 30.200 5.100 30.600 5.500 ;
        RECT 78.200 8.800 78.600 9.200 ;
        RECT 45.400 6.100 45.800 6.500 ;
        RECT 41.400 4.800 41.800 5.200 ;
        RECT 51.800 5.100 52.200 5.500 ;
        RECT 54.200 5.100 54.600 5.500 ;
        RECT 70.200 6.800 70.600 7.200 ;
        RECT 65.400 4.800 65.800 5.200 ;
        RECT 74.200 5.800 74.600 6.200 ;
        RECT 69.400 5.100 69.800 5.500 ;
        RECT 79.000 4.800 79.400 5.200 ;
        RECT 91.000 8.800 91.400 9.200 ;
        RECT 83.800 6.100 84.200 6.500 ;
        RECT 102.200 8.800 102.600 9.200 ;
        RECT 93.400 6.100 93.800 6.500 ;
        RECT 90.200 5.100 90.600 5.500 ;
        RECT 110.200 6.800 110.600 7.200 ;
        RECT 104.600 6.100 105.000 6.500 ;
        RECT 108.600 5.900 109.000 6.300 ;
        RECT 99.800 5.100 100.200 5.500 ;
        RECT 111.000 5.100 111.400 5.500 ;
        RECT 113.400 4.800 113.800 5.200 ;
        RECT 117.400 5.800 117.800 6.200 ;
        RECT 123.000 8.800 123.400 9.200 ;
        RECT 121.400 6.800 121.800 7.200 ;
        RECT 120.600 5.800 121.000 6.200 ;
        RECT 122.200 5.800 122.600 6.200 ;
        RECT 132.600 8.800 133.000 9.200 ;
        RECT 131.000 6.800 131.400 7.200 ;
        RECT 125.400 6.100 125.800 6.500 ;
        RECT 131.800 5.100 132.200 5.500 ;
        RECT 152.600 8.800 153.000 9.200 ;
        RECT 136.600 6.100 137.000 6.500 ;
        RECT 150.200 6.800 150.600 7.200 ;
        RECT 143.000 5.100 143.400 5.500 ;
        RECT 163.000 8.800 163.400 9.200 ;
        RECT 160.600 6.800 161.000 7.200 ;
        RECT 155.000 6.100 155.400 6.500 ;
        RECT 159.000 5.900 159.400 6.300 ;
        RECT 161.400 5.100 161.800 5.500 ;
        RECT 163.800 8.800 164.200 9.200 ;
        RECT 173.400 8.800 173.800 9.200 ;
        RECT 171.800 6.800 172.200 7.200 ;
        RECT 166.200 6.100 166.600 6.500 ;
        RECT 183.000 8.800 183.400 9.200 ;
        RECT 175.800 6.100 176.200 6.500 ;
        RECT 179.800 5.900 180.200 6.300 ;
        RECT 172.600 5.100 173.000 5.500 ;
        RECT 188.600 6.800 189.000 7.200 ;
        RECT 185.400 6.100 185.800 6.500 ;
        RECT 182.200 5.100 182.600 5.500 ;
        RECT 191.800 5.100 192.200 5.500 ;
        RECT 192.600 5.100 193.000 5.500 ;
        RECT 203.000 8.800 203.400 9.200 ;
      LAYER metal2 ;
        RECT 2.200 174.800 2.600 175.200 ;
        RECT 4.600 174.800 5.000 175.200 ;
        RECT 14.200 174.800 14.600 175.200 ;
        RECT 16.600 174.800 17.000 175.200 ;
        RECT 1.400 169.100 1.800 169.200 ;
        RECT 2.200 169.100 2.500 174.800 ;
        RECT 1.400 168.800 2.500 169.100 ;
        RECT 4.600 156.200 4.900 174.800 ;
        RECT 11.000 171.800 11.400 172.200 ;
        RECT 6.200 162.100 6.600 168.900 ;
        RECT 7.000 162.100 7.400 168.900 ;
        RECT 7.800 162.100 8.200 168.900 ;
        RECT 8.600 163.100 9.000 168.900 ;
        RECT 9.400 168.800 9.800 169.200 ;
        RECT 9.400 168.200 9.700 168.800 ;
        RECT 9.400 167.800 9.800 168.200 ;
        RECT 4.600 155.800 5.000 156.200 ;
        RECT 2.200 154.800 2.600 155.200 ;
        RECT 3.800 155.100 4.200 155.200 ;
        RECT 4.600 155.100 5.000 155.200 ;
        RECT 3.800 154.800 5.000 155.100 ;
        RECT 2.200 150.100 2.500 154.800 ;
        RECT 5.400 153.100 5.800 155.900 ;
        RECT 6.200 153.800 6.600 154.200 ;
        RECT 1.400 149.800 2.500 150.100 ;
        RECT 0.600 145.100 1.000 147.900 ;
        RECT 1.400 139.200 1.700 149.800 ;
        RECT 2.200 143.100 2.600 148.900 ;
        RECT 3.000 146.800 3.400 147.200 ;
        RECT 3.800 146.800 4.200 147.200 ;
        RECT 1.400 138.800 1.800 139.200 ;
        RECT 3.000 133.200 3.300 146.800 ;
        RECT 3.800 146.200 4.100 146.800 ;
        RECT 6.200 146.200 6.500 153.800 ;
        RECT 7.000 152.100 7.400 157.900 ;
        RECT 9.400 154.200 9.700 167.800 ;
        RECT 10.200 163.100 10.600 168.900 ;
        RECT 11.000 168.200 11.300 171.800 ;
        RECT 14.200 170.200 14.500 174.800 ;
        RECT 14.200 169.800 14.600 170.200 ;
        RECT 16.600 169.200 16.900 174.800 ;
        RECT 25.400 172.100 25.800 178.900 ;
        RECT 26.200 172.100 26.600 178.900 ;
        RECT 27.000 172.100 27.400 178.900 ;
        RECT 27.800 172.100 28.200 177.900 ;
        RECT 28.600 172.800 29.000 173.200 ;
        RECT 19.000 169.800 19.400 170.200 ;
        RECT 19.000 169.200 19.300 169.800 ;
        RECT 11.000 167.800 11.400 168.200 ;
        RECT 11.000 166.800 11.400 167.200 ;
        RECT 10.200 154.800 10.600 155.200 ;
        RECT 9.400 153.800 9.800 154.200 ;
        RECT 10.200 149.200 10.500 154.800 ;
        RECT 11.000 151.200 11.300 166.800 ;
        RECT 11.800 163.100 12.200 168.900 ;
        RECT 12.600 162.100 13.000 168.900 ;
        RECT 13.400 162.100 13.800 168.900 ;
        RECT 16.600 168.800 17.000 169.200 ;
        RECT 19.000 168.800 19.400 169.200 ;
        RECT 23.000 166.800 23.400 167.200 ;
        RECT 23.000 166.200 23.300 166.800 ;
        RECT 15.800 166.100 16.200 166.200 ;
        RECT 16.600 166.100 17.000 166.200 ;
        RECT 15.800 165.800 17.000 166.100 ;
        RECT 23.000 165.800 23.400 166.200 ;
        RECT 23.800 162.100 24.200 168.900 ;
        RECT 24.600 162.100 25.000 168.900 ;
        RECT 25.400 162.100 25.800 168.900 ;
        RECT 26.200 163.100 26.600 168.900 ;
        RECT 27.000 167.800 27.400 168.200 ;
        RECT 27.000 162.100 27.300 167.800 ;
        RECT 27.800 163.100 28.200 168.900 ;
        RECT 28.600 168.200 28.900 172.800 ;
        RECT 29.400 172.100 29.800 177.900 ;
        RECT 30.200 173.800 30.600 174.200 ;
        RECT 30.200 170.200 30.500 173.800 ;
        RECT 31.000 172.100 31.400 177.900 ;
        RECT 31.800 172.100 32.200 178.900 ;
        RECT 32.600 172.100 33.000 178.900 ;
        RECT 33.400 174.800 33.800 175.200 ;
        RECT 35.000 174.800 35.400 175.200 ;
        RECT 37.400 174.800 37.800 175.200 ;
        RECT 39.800 174.800 40.200 175.200 ;
        RECT 49.400 174.800 49.800 175.200 ;
        RECT 30.200 169.800 30.600 170.200 ;
        RECT 28.600 167.800 29.000 168.200 ;
        RECT 28.600 166.800 29.000 167.200 ;
        RECT 28.600 164.200 28.900 166.800 ;
        RECT 28.600 163.800 29.000 164.200 ;
        RECT 29.400 163.100 29.800 168.900 ;
        RECT 30.200 162.100 30.600 168.900 ;
        RECT 31.000 162.100 31.400 168.900 ;
        RECT 33.400 166.200 33.700 174.800 ;
        RECT 35.000 174.200 35.300 174.800 ;
        RECT 37.400 174.200 37.700 174.800 ;
        RECT 35.000 173.800 35.400 174.200 ;
        RECT 37.400 173.800 37.800 174.200 ;
        RECT 35.800 169.100 36.200 169.200 ;
        RECT 36.600 169.100 37.000 169.200 ;
        RECT 35.800 168.800 37.000 169.100 ;
        RECT 39.800 167.200 40.100 174.800 ;
        RECT 44.600 171.800 45.000 172.200 ;
        RECT 39.800 166.800 40.200 167.200 ;
        RECT 33.400 165.800 33.800 166.200 ;
        RECT 26.200 161.800 27.300 162.100 ;
        RECT 11.800 152.100 12.200 157.900 ;
        RECT 16.600 154.800 17.000 155.200 ;
        RECT 17.400 155.100 17.800 155.200 ;
        RECT 18.100 155.100 18.500 155.200 ;
        RECT 17.400 154.800 18.500 155.100 ;
        RECT 21.400 154.800 21.800 155.200 ;
        RECT 16.600 153.200 16.900 154.800 ;
        RECT 13.400 152.800 13.800 153.200 ;
        RECT 15.000 152.800 15.400 153.200 ;
        RECT 16.600 152.800 17.000 153.200 ;
        RECT 11.000 150.800 11.400 151.200 ;
        RECT 3.800 145.800 4.200 146.200 ;
        RECT 6.200 145.800 6.600 146.200 ;
        RECT 7.000 143.100 7.400 148.900 ;
        RECT 9.400 148.800 9.800 149.200 ;
        RECT 10.200 148.800 10.600 149.200 ;
        RECT 9.400 148.200 9.700 148.800 ;
        RECT 9.400 147.800 9.800 148.200 ;
        RECT 13.400 147.200 13.700 152.800 ;
        RECT 15.000 150.200 15.300 152.800 ;
        RECT 15.800 151.800 16.200 152.200 ;
        RECT 15.000 149.800 15.400 150.200 ;
        RECT 14.200 149.100 14.600 149.200 ;
        RECT 15.000 149.100 15.400 149.200 ;
        RECT 14.200 148.800 15.400 149.100 ;
        RECT 15.800 148.200 16.100 151.800 ;
        RECT 15.800 147.800 16.200 148.200 ;
        RECT 16.600 147.800 17.000 148.200 ;
        RECT 16.600 147.200 16.900 147.800 ;
        RECT 21.400 147.200 21.700 154.800 ;
        RECT 23.000 152.100 23.400 158.900 ;
        RECT 23.800 152.100 24.200 158.900 ;
        RECT 24.600 152.100 25.000 158.900 ;
        RECT 25.400 152.100 25.800 157.900 ;
        RECT 26.200 153.200 26.500 161.800 ;
        RECT 26.200 152.800 26.600 153.200 ;
        RECT 10.200 146.800 10.600 147.200 ;
        RECT 11.000 147.100 11.400 147.200 ;
        RECT 11.800 147.100 12.200 147.200 ;
        RECT 11.000 146.800 12.200 147.100 ;
        RECT 12.600 146.800 13.000 147.200 ;
        RECT 13.400 146.800 13.800 147.200 ;
        RECT 16.600 146.800 17.000 147.200 ;
        RECT 17.400 147.100 17.800 147.200 ;
        RECT 18.200 147.100 18.600 147.200 ;
        RECT 17.400 146.800 18.600 147.100 ;
        RECT 19.000 147.100 19.400 147.200 ;
        RECT 19.800 147.100 20.200 147.200 ;
        RECT 19.000 146.800 20.200 147.100 ;
        RECT 21.400 146.800 21.800 147.200 ;
        RECT 10.200 144.200 10.500 146.800 ;
        RECT 11.000 146.100 11.400 146.200 ;
        RECT 11.800 146.100 12.200 146.200 ;
        RECT 11.000 145.800 12.200 146.100 ;
        RECT 12.600 145.200 12.900 146.800 ;
        RECT 13.400 145.800 13.800 146.200 ;
        RECT 14.200 145.800 14.600 146.200 ;
        RECT 18.200 145.800 18.600 146.200 ;
        RECT 20.600 145.800 21.000 146.200 ;
        RECT 13.400 145.200 13.700 145.800 ;
        RECT 12.600 144.800 13.000 145.200 ;
        RECT 13.400 144.800 13.800 145.200 ;
        RECT 10.200 143.800 10.600 144.200 ;
        RECT 3.000 132.800 3.400 133.200 ;
        RECT 0.600 125.100 1.000 127.900 ;
        RECT 2.200 123.100 2.600 128.900 ;
        RECT 3.000 128.200 3.300 132.800 ;
        RECT 6.200 132.100 6.600 138.900 ;
        RECT 7.000 132.100 7.400 138.900 ;
        RECT 7.800 132.100 8.200 138.900 ;
        RECT 8.600 132.100 9.000 137.900 ;
        RECT 9.400 133.800 9.800 134.200 ;
        RECT 9.400 133.200 9.700 133.800 ;
        RECT 9.400 132.800 9.800 133.200 ;
        RECT 10.200 132.100 10.600 137.900 ;
        RECT 11.000 133.800 11.400 134.200 ;
        RECT 11.000 131.200 11.300 133.800 ;
        RECT 11.800 132.100 12.200 137.900 ;
        RECT 12.600 132.100 13.000 138.900 ;
        RECT 13.400 132.100 13.800 138.900 ;
        RECT 11.000 130.800 11.400 131.200 ;
        RECT 3.000 127.800 3.400 128.200 ;
        RECT 0.600 113.100 1.000 115.900 ;
        RECT 2.200 112.100 2.600 117.900 ;
        RECT 3.000 114.200 3.300 127.800 ;
        RECT 5.400 126.800 5.800 127.200 ;
        RECT 5.400 126.200 5.700 126.800 ;
        RECT 5.400 125.800 5.800 126.200 ;
        RECT 7.000 123.100 7.400 128.900 ;
        RECT 11.000 128.800 11.400 129.200 ;
        RECT 11.000 128.200 11.300 128.800 ;
        RECT 11.000 127.800 11.400 128.200 ;
        RECT 11.800 127.100 12.200 127.200 ;
        RECT 12.600 127.100 13.000 127.200 ;
        RECT 11.800 126.800 13.000 127.100 ;
        RECT 12.600 126.100 13.000 126.200 ;
        RECT 13.400 126.100 13.800 126.200 ;
        RECT 12.600 125.800 13.800 126.100 ;
        RECT 5.400 114.800 5.800 115.200 ;
        RECT 3.000 113.800 3.400 114.200 ;
        RECT 5.400 109.200 5.700 114.800 ;
        RECT 7.000 112.100 7.400 117.900 ;
        RECT 10.200 113.100 10.600 115.900 ;
        RECT 11.000 114.800 11.400 115.200 ;
        RECT 11.000 114.200 11.300 114.800 ;
        RECT 11.000 113.800 11.400 114.200 ;
        RECT 9.400 111.800 9.800 112.200 ;
        RECT 11.800 112.100 12.200 117.900 ;
        RECT 0.600 108.800 1.000 109.200 ;
        RECT 0.600 108.200 0.900 108.800 ;
        RECT 0.600 107.800 1.000 108.200 ;
        RECT 3.000 103.100 3.400 108.900 ;
        RECT 5.400 108.800 5.800 109.200 ;
        RECT 9.400 109.100 9.700 111.800 ;
        RECT 6.200 106.800 6.600 107.200 ;
        RECT 6.200 99.200 6.500 106.800 ;
        RECT 7.000 105.900 7.400 106.300 ;
        RECT 7.000 105.200 7.300 105.900 ;
        RECT 7.000 104.800 7.400 105.200 ;
        RECT 7.800 103.100 8.200 108.900 ;
        RECT 9.400 108.800 10.500 109.100 ;
        RECT 10.200 108.200 10.500 108.800 ;
        RECT 9.400 105.100 9.800 107.900 ;
        RECT 10.200 107.800 10.600 108.200 ;
        RECT 12.600 107.200 12.900 125.800 ;
        RECT 14.200 116.100 14.500 145.800 ;
        RECT 18.200 145.200 18.500 145.800 ;
        RECT 18.200 144.800 18.600 145.200 ;
        RECT 19.000 144.800 19.400 145.200 ;
        RECT 19.000 139.200 19.300 144.800 ;
        RECT 20.600 144.200 20.900 145.800 ;
        RECT 21.400 145.200 21.700 146.800 ;
        RECT 21.400 144.800 21.800 145.200 ;
        RECT 22.200 145.100 22.600 147.900 ;
        RECT 23.000 146.800 23.400 147.200 ;
        RECT 20.600 143.800 21.000 144.200 ;
        RECT 19.800 141.800 20.200 142.200 ;
        RECT 19.000 138.800 19.400 139.200 ;
        RECT 18.200 135.800 18.600 136.200 ;
        RECT 18.200 135.200 18.500 135.800 ;
        RECT 15.800 134.800 16.200 135.200 ;
        RECT 18.200 134.800 18.600 135.200 ;
        RECT 15.800 134.200 16.100 134.800 ;
        RECT 19.800 134.200 20.100 141.800 ;
        RECT 20.600 139.100 21.000 139.200 ;
        RECT 21.400 139.100 21.800 139.200 ;
        RECT 20.600 138.800 21.800 139.100 ;
        RECT 15.800 133.800 16.200 134.200 ;
        RECT 19.800 133.800 20.200 134.200 ;
        RECT 15.000 129.800 15.400 130.200 ;
        RECT 15.000 128.200 15.300 129.800 ;
        RECT 15.000 127.800 15.400 128.200 ;
        RECT 15.000 126.200 15.300 127.800 ;
        RECT 15.000 125.800 15.400 126.200 ;
        RECT 15.800 125.800 16.200 126.200 ;
        RECT 15.800 125.200 16.100 125.800 ;
        RECT 15.800 124.800 16.200 125.200 ;
        RECT 16.600 125.100 17.000 127.900 ;
        RECT 17.400 126.800 17.800 127.200 ;
        RECT 14.200 115.800 15.300 116.100 ;
        RECT 14.200 114.800 14.600 115.200 ;
        RECT 14.200 113.200 14.500 114.800 ;
        RECT 14.200 112.800 14.600 113.200 ;
        RECT 11.800 107.100 12.200 107.200 ;
        RECT 12.600 107.100 13.000 107.200 ;
        RECT 11.800 106.800 13.000 107.100 ;
        RECT 15.000 106.200 15.300 115.800 ;
        RECT 16.600 112.100 17.000 117.900 ;
        RECT 17.400 117.200 17.700 126.800 ;
        RECT 18.200 123.100 18.600 128.900 ;
        RECT 19.800 128.200 20.100 133.800 ;
        RECT 23.000 133.200 23.300 146.800 ;
        RECT 23.800 143.100 24.200 148.900 ;
        RECT 26.200 148.200 26.500 152.800 ;
        RECT 27.000 152.100 27.400 157.900 ;
        RECT 27.800 153.800 28.200 154.200 ;
        RECT 27.800 149.200 28.100 153.800 ;
        RECT 28.600 152.100 29.000 157.900 ;
        RECT 29.400 152.100 29.800 158.900 ;
        RECT 30.200 152.100 30.600 158.900 ;
        RECT 33.400 155.200 33.700 165.800 ;
        RECT 35.000 164.800 35.400 165.200 ;
        RECT 35.000 155.200 35.300 164.800 ;
        RECT 41.400 162.100 41.800 168.900 ;
        RECT 42.200 162.100 42.600 168.900 ;
        RECT 43.000 162.100 43.400 168.900 ;
        RECT 43.800 163.100 44.200 168.900 ;
        RECT 44.600 168.200 44.900 171.800 ;
        RECT 49.400 171.200 49.700 174.800 ;
        RECT 50.200 172.100 50.600 178.900 ;
        RECT 51.000 172.100 51.400 178.900 ;
        RECT 51.800 172.100 52.200 178.900 ;
        RECT 52.600 172.100 53.000 177.900 ;
        RECT 53.400 172.800 53.800 173.200 ;
        RECT 53.400 172.200 53.700 172.800 ;
        RECT 53.400 171.800 53.800 172.200 ;
        RECT 54.200 172.100 54.600 177.900 ;
        RECT 55.000 173.800 55.400 174.200 ;
        RECT 49.400 170.800 49.800 171.200 ;
        RECT 51.000 170.800 51.400 171.200 ;
        RECT 44.600 167.800 45.000 168.200 ;
        RECT 33.400 154.800 33.800 155.200 ;
        RECT 35.000 154.800 35.400 155.200 ;
        RECT 38.200 154.800 38.600 155.200 ;
        RECT 33.400 150.100 33.700 154.800 ;
        RECT 33.400 149.800 34.500 150.100 ;
        RECT 27.800 148.800 28.200 149.200 ;
        RECT 26.200 147.800 26.600 148.200 ;
        RECT 24.600 146.800 25.000 147.200 ;
        RECT 24.600 146.300 24.900 146.800 ;
        RECT 24.600 145.900 25.000 146.300 ;
        RECT 28.600 143.100 29.000 148.900 ;
        RECT 31.800 145.100 32.200 147.900 ;
        RECT 33.400 143.100 33.800 148.900 ;
        RECT 30.200 142.100 30.600 142.200 ;
        RECT 31.000 142.100 31.400 142.200 ;
        RECT 30.200 141.800 31.400 142.100 ;
        RECT 25.400 134.800 25.800 135.200 ;
        RECT 25.400 134.200 25.700 134.800 ;
        RECT 25.400 133.800 25.800 134.200 ;
        RECT 23.000 132.800 23.400 133.200 ;
        RECT 26.200 132.100 26.600 138.900 ;
        RECT 27.000 132.100 27.400 138.900 ;
        RECT 27.800 132.100 28.200 138.900 ;
        RECT 28.600 132.100 29.000 137.900 ;
        RECT 29.400 132.800 29.800 133.200 ;
        RECT 29.400 132.200 29.700 132.800 ;
        RECT 29.400 131.800 29.800 132.200 ;
        RECT 30.200 132.100 30.600 137.900 ;
        RECT 31.000 133.800 31.400 134.200 ;
        RECT 19.800 127.800 20.200 128.200 ;
        RECT 19.800 125.800 20.200 126.200 ;
        RECT 21.400 125.800 21.800 126.200 ;
        RECT 19.800 125.200 20.100 125.800 ;
        RECT 19.800 124.800 20.200 125.200 ;
        RECT 17.400 116.800 17.800 117.200 ;
        RECT 21.400 115.200 21.700 125.800 ;
        RECT 23.000 123.100 23.400 128.900 ;
        RECT 25.400 128.800 25.800 129.200 ;
        RECT 27.000 128.800 27.400 129.200 ;
        RECT 29.400 128.800 29.800 129.200 ;
        RECT 25.400 127.200 25.700 128.800 ;
        RECT 25.400 126.800 25.800 127.200 ;
        RECT 26.200 126.800 26.600 127.200 ;
        RECT 26.200 126.200 26.500 126.800 ;
        RECT 27.000 126.200 27.300 128.800 ;
        RECT 28.600 127.800 29.000 128.200 ;
        RECT 24.600 125.800 25.000 126.200 ;
        RECT 26.200 125.800 26.600 126.200 ;
        RECT 27.000 125.800 27.400 126.200 ;
        RECT 22.200 115.800 22.600 116.200 ;
        RECT 22.200 115.200 22.500 115.800 ;
        RECT 24.600 115.200 24.900 125.800 ;
        RECT 27.000 125.100 27.400 125.200 ;
        RECT 27.800 125.100 28.200 125.200 ;
        RECT 27.000 124.800 28.200 125.100 ;
        RECT 19.800 115.100 20.200 115.200 ;
        RECT 20.600 115.100 21.000 115.200 ;
        RECT 19.800 114.800 21.000 115.100 ;
        RECT 21.400 114.800 21.800 115.200 ;
        RECT 22.200 114.800 22.600 115.200 ;
        RECT 24.600 114.800 25.000 115.200 ;
        RECT 16.600 109.800 17.000 110.200 ;
        RECT 16.600 106.200 16.900 109.800 ;
        RECT 18.200 109.100 18.600 109.200 ;
        RECT 19.000 109.100 19.400 109.200 ;
        RECT 18.200 108.800 19.400 109.100 ;
        RECT 17.400 107.800 17.800 108.200 ;
        RECT 17.400 107.200 17.700 107.800 ;
        RECT 17.400 106.800 17.800 107.200 ;
        RECT 21.400 106.200 21.700 114.800 ;
        RECT 23.000 113.100 23.400 113.200 ;
        RECT 23.800 113.100 24.200 113.200 ;
        RECT 26.200 113.100 26.600 115.900 ;
        RECT 27.000 114.800 27.400 115.200 ;
        RECT 27.000 114.200 27.300 114.800 ;
        RECT 27.000 113.800 27.400 114.200 ;
        RECT 23.000 112.800 24.200 113.100 ;
        RECT 27.800 112.100 28.200 117.900 ;
        RECT 22.200 108.800 22.600 109.200 ;
        RECT 27.800 108.800 28.200 109.200 ;
        RECT 22.200 108.200 22.500 108.800 ;
        RECT 27.800 108.200 28.100 108.800 ;
        RECT 22.200 107.800 22.600 108.200 ;
        RECT 26.200 108.100 26.600 108.200 ;
        RECT 27.000 108.100 27.400 108.200 ;
        RECT 26.200 107.800 27.400 108.100 ;
        RECT 27.800 107.800 28.200 108.200 ;
        RECT 23.800 107.100 24.200 107.200 ;
        RECT 24.600 107.100 25.000 107.200 ;
        RECT 23.800 106.800 25.000 107.100 ;
        RECT 12.600 106.100 13.000 106.200 ;
        RECT 13.400 106.100 13.800 106.200 ;
        RECT 12.600 105.800 13.800 106.100 ;
        RECT 15.000 105.800 15.400 106.200 ;
        RECT 16.600 105.800 17.000 106.200 ;
        RECT 17.400 105.800 17.800 106.200 ;
        RECT 20.600 105.800 21.000 106.200 ;
        RECT 21.400 105.800 21.800 106.200 ;
        RECT 15.000 105.200 15.300 105.800 ;
        RECT 12.600 104.800 13.000 105.200 ;
        RECT 15.000 104.800 15.400 105.200 ;
        RECT 12.600 104.200 12.900 104.800 ;
        RECT 11.000 103.800 11.400 104.200 ;
        RECT 12.600 103.800 13.000 104.200 ;
        RECT 11.000 103.200 11.300 103.800 ;
        RECT 11.000 102.800 11.400 103.200 ;
        RECT 6.200 98.800 6.600 99.200 ;
        RECT 7.800 93.100 8.200 95.900 ;
        RECT 8.600 93.800 9.000 94.200 ;
        RECT 6.200 91.800 6.600 92.200 ;
        RECT 0.600 88.800 1.000 89.200 ;
        RECT 0.600 88.200 0.900 88.800 ;
        RECT 0.600 87.800 1.000 88.200 ;
        RECT 3.000 83.100 3.400 88.900 ;
        RECT 6.200 87.200 6.500 91.800 ;
        RECT 6.200 86.800 6.600 87.200 ;
        RECT 7.000 86.800 7.400 87.200 ;
        RECT 7.000 86.300 7.300 86.800 ;
        RECT 7.000 85.900 7.400 86.300 ;
        RECT 7.800 83.100 8.200 88.900 ;
        RECT 8.600 87.200 8.900 93.800 ;
        RECT 9.400 92.100 9.800 97.900 ;
        RECT 11.800 95.100 12.200 95.200 ;
        RECT 12.600 95.100 13.000 95.200 ;
        RECT 11.800 94.800 13.000 95.100 ;
        RECT 14.200 92.100 14.600 97.900 ;
        RECT 15.000 90.200 15.300 104.800 ;
        RECT 17.400 94.200 17.700 105.800 ;
        RECT 20.600 103.200 20.900 105.800 ;
        RECT 21.400 105.200 21.700 105.800 ;
        RECT 21.400 104.800 21.800 105.200 ;
        RECT 20.600 102.800 21.000 103.200 ;
        RECT 18.200 95.800 18.600 96.200 ;
        RECT 22.200 96.100 22.600 96.200 ;
        RECT 23.000 96.100 23.400 96.200 ;
        RECT 22.200 95.800 23.400 96.100 ;
        RECT 18.200 95.200 18.500 95.800 ;
        RECT 18.200 94.800 18.600 95.200 ;
        RECT 19.000 95.100 19.400 95.200 ;
        RECT 19.800 95.100 20.200 95.200 ;
        RECT 19.000 94.800 20.200 95.100 ;
        RECT 20.600 94.800 21.000 95.200 ;
        RECT 22.200 94.800 22.600 95.200 ;
        RECT 20.600 94.200 20.900 94.800 ;
        RECT 15.800 94.100 16.200 94.200 ;
        RECT 16.600 94.100 17.000 94.200 ;
        RECT 15.800 93.800 17.000 94.100 ;
        RECT 17.400 93.800 17.800 94.200 ;
        RECT 20.600 93.800 21.000 94.200 ;
        RECT 15.000 89.800 15.400 90.200 ;
        RECT 17.400 89.200 17.700 93.800 ;
        RECT 20.600 91.800 21.000 92.200 ;
        RECT 19.800 89.800 20.200 90.200 ;
        RECT 15.000 88.800 15.400 89.200 ;
        RECT 17.400 88.800 17.800 89.200 ;
        RECT 8.600 86.800 9.000 87.200 ;
        RECT 9.400 85.100 9.800 87.900 ;
        RECT 10.200 87.800 10.600 88.200 ;
        RECT 10.200 87.200 10.500 87.800 ;
        RECT 10.200 86.800 10.600 87.200 ;
        RECT 11.800 86.800 12.200 87.200 ;
        RECT 11.800 86.200 12.100 86.800 ;
        RECT 11.800 85.800 12.200 86.200 ;
        RECT 14.200 85.800 14.600 86.200 ;
        RECT 11.800 84.800 12.200 85.200 ;
        RECT 9.400 81.800 9.800 82.200 ;
        RECT 9.400 79.200 9.700 81.800 ;
        RECT 11.800 81.200 12.100 84.800 ;
        RECT 14.200 81.200 14.500 85.800 ;
        RECT 11.800 80.800 12.200 81.200 ;
        RECT 14.200 80.800 14.600 81.200 ;
        RECT 9.400 78.800 9.800 79.200 ;
        RECT 0.600 73.100 1.000 75.900 ;
        RECT 2.200 72.100 2.600 77.900 ;
        RECT 4.600 75.100 5.000 75.200 ;
        RECT 5.400 75.100 5.800 75.200 ;
        RECT 4.600 74.800 5.800 75.100 ;
        RECT 3.000 72.800 3.400 73.200 ;
        RECT 0.600 65.100 1.000 67.900 ;
        RECT 2.200 63.100 2.600 68.900 ;
        RECT 3.000 68.200 3.300 72.800 ;
        RECT 7.000 72.100 7.400 77.900 ;
        RECT 15.000 75.200 15.300 88.800 ;
        RECT 18.200 87.800 18.600 88.200 ;
        RECT 19.000 87.800 19.400 88.200 ;
        RECT 15.800 86.800 16.200 87.200 ;
        RECT 17.400 86.800 17.800 87.200 ;
        RECT 15.800 86.200 16.100 86.800 ;
        RECT 17.400 86.200 17.700 86.800 ;
        RECT 18.200 86.200 18.500 87.800 ;
        RECT 19.000 87.200 19.300 87.800 ;
        RECT 19.000 86.800 19.400 87.200 ;
        RECT 15.800 85.800 16.200 86.200 ;
        RECT 17.400 85.800 17.800 86.200 ;
        RECT 18.200 85.800 18.600 86.200 ;
        RECT 15.800 84.800 16.200 85.200 ;
        RECT 15.800 83.200 16.100 84.800 ;
        RECT 15.800 82.800 16.200 83.200 ;
        RECT 18.200 82.800 18.600 83.200 ;
        RECT 16.600 81.800 17.000 82.200 ;
        RECT 15.800 76.100 16.200 76.200 ;
        RECT 16.600 76.100 16.900 81.800 ;
        RECT 15.800 75.800 16.900 76.100 ;
        RECT 18.200 75.200 18.500 82.800 ;
        RECT 11.800 74.800 12.200 75.200 ;
        RECT 12.600 75.100 13.000 75.200 ;
        RECT 13.400 75.100 13.800 75.200 ;
        RECT 12.600 74.800 13.800 75.100 ;
        RECT 14.200 74.800 14.600 75.200 ;
        RECT 15.000 74.800 15.400 75.200 ;
        RECT 15.800 75.100 16.200 75.200 ;
        RECT 16.600 75.100 17.000 75.200 ;
        RECT 15.800 74.800 17.000 75.100 ;
        RECT 18.200 74.800 18.600 75.200 ;
        RECT 11.800 74.200 12.100 74.800 ;
        RECT 14.200 74.200 14.500 74.800 ;
        RECT 11.800 73.800 12.200 74.200 ;
        RECT 14.200 73.800 14.600 74.200 ;
        RECT 15.000 71.200 15.300 74.800 ;
        RECT 18.200 73.800 18.600 74.200 ;
        RECT 18.200 73.200 18.500 73.800 ;
        RECT 18.200 72.800 18.600 73.200 ;
        RECT 19.000 73.100 19.400 75.900 ;
        RECT 15.000 70.800 15.400 71.200 ;
        RECT 9.400 69.100 9.800 69.200 ;
        RECT 10.200 69.100 10.600 69.200 ;
        RECT 3.000 67.800 3.400 68.200 ;
        RECT 4.600 66.100 5.000 66.200 ;
        RECT 5.400 66.100 5.800 66.200 ;
        RECT 4.600 65.800 5.800 66.100 ;
        RECT 6.200 65.800 6.600 66.200 ;
        RECT 6.200 65.200 6.500 65.800 ;
        RECT 6.200 64.800 6.600 65.200 ;
        RECT 0.600 53.100 1.000 55.900 ;
        RECT 2.200 52.100 2.600 57.900 ;
        RECT 3.800 54.800 4.200 55.200 ;
        RECT 3.000 53.800 3.400 54.200 ;
        RECT 3.000 53.200 3.300 53.800 ;
        RECT 3.000 52.800 3.400 53.200 ;
        RECT 0.600 35.100 1.000 35.200 ;
        RECT 1.400 35.100 1.800 35.200 ;
        RECT 0.600 34.800 1.800 35.100 ;
        RECT 0.600 32.800 1.000 33.200 ;
        RECT 2.200 33.100 2.600 35.900 ;
        RECT 3.000 34.200 3.300 52.800 ;
        RECT 3.800 51.200 4.100 54.800 ;
        RECT 3.800 50.800 4.200 51.200 ;
        RECT 6.200 49.200 6.500 64.800 ;
        RECT 7.000 63.100 7.400 68.900 ;
        RECT 9.400 68.800 10.600 69.100 ;
        RECT 15.000 68.800 15.400 69.200 ;
        RECT 15.000 67.200 15.300 68.800 ;
        RECT 10.200 66.800 10.600 67.200 ;
        RECT 12.600 66.800 13.000 67.200 ;
        RECT 13.400 67.100 13.800 67.200 ;
        RECT 14.200 67.100 14.600 67.200 ;
        RECT 13.400 66.800 14.600 67.100 ;
        RECT 15.000 66.800 15.400 67.200 ;
        RECT 10.200 65.200 10.500 66.800 ;
        RECT 11.000 66.100 11.400 66.200 ;
        RECT 11.800 66.100 12.200 66.200 ;
        RECT 11.000 65.800 12.200 66.100 ;
        RECT 10.200 64.800 10.600 65.200 ;
        RECT 12.600 64.100 12.900 66.800 ;
        RECT 13.400 65.800 13.800 66.200 ;
        RECT 15.000 65.800 15.400 66.200 ;
        RECT 13.400 65.200 13.700 65.800 ;
        RECT 13.400 64.800 13.800 65.200 ;
        RECT 12.600 63.800 13.700 64.100 ;
        RECT 9.400 60.800 9.800 61.200 ;
        RECT 9.400 59.200 9.700 60.800 ;
        RECT 9.400 58.800 9.800 59.200 ;
        RECT 12.600 58.800 13.000 59.200 ;
        RECT 7.000 52.100 7.400 57.900 ;
        RECT 10.200 53.100 10.600 55.900 ;
        RECT 11.000 53.800 11.400 54.200 ;
        RECT 11.000 53.200 11.300 53.800 ;
        RECT 11.000 52.800 11.400 53.200 ;
        RECT 7.800 51.800 8.200 52.200 ;
        RECT 8.600 52.100 9.000 52.200 ;
        RECT 9.400 52.100 9.800 52.200 ;
        RECT 11.800 52.100 12.200 57.900 ;
        RECT 8.600 51.800 9.800 52.100 ;
        RECT 6.200 48.800 6.600 49.200 ;
        RECT 7.800 48.200 8.100 51.800 ;
        RECT 11.000 50.800 11.400 51.200 ;
        RECT 11.000 49.200 11.300 50.800 ;
        RECT 11.000 48.800 11.400 49.200 ;
        RECT 7.800 47.800 8.200 48.200 ;
        RECT 12.600 47.200 12.900 58.800 ;
        RECT 13.400 54.200 13.700 63.800 ;
        RECT 14.200 56.800 14.600 57.200 ;
        RECT 14.200 55.200 14.500 56.800 ;
        RECT 14.200 54.800 14.600 55.200 ;
        RECT 13.400 53.800 13.800 54.200 ;
        RECT 9.400 46.800 9.800 47.200 ;
        RECT 12.600 46.800 13.000 47.200 ;
        RECT 13.400 46.800 13.800 47.200 ;
        RECT 9.400 46.200 9.700 46.800 ;
        RECT 9.400 45.800 9.800 46.200 ;
        RECT 11.800 46.100 12.200 46.200 ;
        RECT 12.600 46.100 13.000 46.200 ;
        RECT 11.800 45.800 13.000 46.100 ;
        RECT 11.000 39.100 11.400 39.200 ;
        RECT 11.800 39.100 12.200 39.200 ;
        RECT 11.000 38.800 12.200 39.100 ;
        RECT 3.000 33.800 3.400 34.200 ;
        RECT 0.600 29.200 0.900 32.800 ;
        RECT 3.800 32.100 4.200 37.900 ;
        RECT 5.400 36.800 5.800 37.200 ;
        RECT 5.400 35.200 5.700 36.800 ;
        RECT 5.400 34.800 5.800 35.200 ;
        RECT 6.200 33.800 6.600 34.200 ;
        RECT 0.600 28.800 1.000 29.200 ;
        RECT 3.000 23.100 3.400 28.900 ;
        RECT 6.200 27.200 6.500 33.800 ;
        RECT 7.000 31.800 7.400 32.200 ;
        RECT 8.600 32.100 9.000 37.900 ;
        RECT 12.600 35.200 12.900 45.800 ;
        RECT 13.400 39.200 13.700 46.800 ;
        RECT 15.000 46.200 15.300 65.800 ;
        RECT 15.800 65.100 16.200 67.900 ;
        RECT 16.600 66.800 17.000 67.200 ;
        RECT 16.600 65.200 16.900 66.800 ;
        RECT 16.600 64.800 17.000 65.200 ;
        RECT 17.400 63.100 17.800 68.900 ;
        RECT 18.200 66.200 18.500 72.800 ;
        RECT 19.000 67.800 19.400 68.200 ;
        RECT 19.000 66.200 19.300 67.800 ;
        RECT 18.200 65.800 18.600 66.200 ;
        RECT 19.000 65.800 19.400 66.200 ;
        RECT 16.600 52.100 17.000 57.900 ;
        RECT 19.000 56.800 19.400 57.200 ;
        RECT 18.200 55.800 18.600 56.200 ;
        RECT 15.800 46.800 16.200 47.200 ;
        RECT 15.000 45.800 15.400 46.200 ;
        RECT 15.000 45.200 15.300 45.800 ;
        RECT 15.000 44.800 15.400 45.200 ;
        RECT 13.400 38.800 13.800 39.200 ;
        RECT 15.800 37.200 16.100 46.800 ;
        RECT 18.200 46.200 18.500 55.800 ;
        RECT 19.000 55.200 19.300 56.800 ;
        RECT 19.800 56.200 20.100 89.800 ;
        RECT 20.600 88.200 20.900 91.800 ;
        RECT 21.400 90.800 21.800 91.200 ;
        RECT 21.400 89.200 21.700 90.800 ;
        RECT 21.400 88.800 21.800 89.200 ;
        RECT 20.600 87.800 21.000 88.200 ;
        RECT 22.200 86.200 22.500 94.800 ;
        RECT 23.800 94.200 24.100 106.800 ;
        RECT 28.600 106.200 28.900 127.800 ;
        RECT 29.400 125.200 29.700 128.800 ;
        RECT 31.000 128.200 31.300 133.800 ;
        RECT 31.800 132.100 32.200 137.900 ;
        RECT 32.600 132.100 33.000 138.900 ;
        RECT 33.400 132.100 33.800 138.900 ;
        RECT 34.200 135.200 34.500 149.800 ;
        RECT 34.200 134.800 34.600 135.200 ;
        RECT 31.000 127.800 31.400 128.200 ;
        RECT 31.000 126.800 31.400 127.200 ;
        RECT 31.000 126.200 31.300 126.800 ;
        RECT 31.000 125.800 31.400 126.200 ;
        RECT 29.400 124.800 29.800 125.200 ;
        RECT 31.800 125.100 32.200 127.900 ;
        RECT 33.400 123.100 33.800 128.900 ;
        RECT 35.000 126.200 35.300 154.800 ;
        RECT 35.800 153.800 36.200 154.200 ;
        RECT 35.800 153.200 36.100 153.800 ;
        RECT 38.200 153.200 38.500 154.800 ;
        RECT 35.800 152.800 36.200 153.200 ;
        RECT 38.200 152.800 38.600 153.200 ;
        RECT 39.800 152.800 40.200 153.200 ;
        RECT 40.600 153.100 41.000 155.900 ;
        RECT 36.600 151.800 37.000 152.200 ;
        RECT 35.800 147.800 36.200 148.200 ;
        RECT 35.800 147.200 36.100 147.800 ;
        RECT 35.800 146.800 36.200 147.200 ;
        RECT 36.600 146.200 36.900 151.800 ;
        RECT 36.600 145.800 37.000 146.200 ;
        RECT 38.200 143.100 38.600 148.900 ;
        RECT 39.800 147.200 40.100 152.800 ;
        RECT 42.200 152.100 42.600 157.900 ;
        RECT 43.800 155.800 44.200 156.200 ;
        RECT 43.800 155.200 44.100 155.800 ;
        RECT 43.800 154.800 44.200 155.200 ;
        RECT 44.600 154.200 44.900 167.800 ;
        RECT 45.400 163.100 45.800 168.900 ;
        RECT 46.200 166.800 46.600 167.200 ;
        RECT 46.200 163.200 46.500 166.800 ;
        RECT 46.200 162.800 46.600 163.200 ;
        RECT 47.000 163.100 47.400 168.900 ;
        RECT 47.800 162.100 48.200 168.900 ;
        RECT 48.600 162.100 49.000 168.900 ;
        RECT 51.000 166.200 51.300 170.800 ;
        RECT 53.400 166.800 53.800 167.200 ;
        RECT 53.400 166.200 53.700 166.800 ;
        RECT 51.000 166.100 51.400 166.200 ;
        RECT 51.800 166.100 52.200 166.200 ;
        RECT 51.000 165.800 52.200 166.100 ;
        RECT 53.400 165.800 53.800 166.200 ;
        RECT 55.000 160.200 55.300 173.800 ;
        RECT 55.800 172.100 56.200 177.900 ;
        RECT 56.600 172.100 57.000 178.900 ;
        RECT 57.400 172.100 57.800 178.900 ;
        RECT 60.600 174.800 61.000 175.200 ;
        RECT 57.400 170.800 57.800 171.200 ;
        RECT 57.400 167.200 57.700 170.800 ;
        RECT 60.600 169.200 60.900 174.800 ;
        RECT 62.200 172.100 62.600 172.200 ;
        RECT 64.600 172.100 65.000 177.900 ;
        RECT 67.000 175.100 67.400 175.200 ;
        RECT 67.800 175.100 68.200 175.200 ;
        RECT 67.000 174.800 68.200 175.100 ;
        RECT 65.400 173.800 65.800 174.200 ;
        RECT 66.200 173.800 66.600 174.200 ;
        RECT 62.200 171.800 63.300 172.100 ;
        RECT 60.600 168.800 61.000 169.200 ;
        RECT 63.000 167.200 63.300 171.800 ;
        RECT 65.400 169.200 65.700 173.800 ;
        RECT 66.200 173.200 66.500 173.800 ;
        RECT 66.200 172.800 66.600 173.200 ;
        RECT 65.400 168.800 65.800 169.200 ;
        RECT 57.400 166.800 57.800 167.200 ;
        RECT 58.200 166.800 58.600 167.200 ;
        RECT 63.000 166.800 63.400 167.200 ;
        RECT 64.600 166.800 65.000 167.200 ;
        RECT 57.400 166.200 57.700 166.800 ;
        RECT 57.400 165.800 57.800 166.200 ;
        RECT 58.200 165.200 58.500 166.800 ;
        RECT 59.000 165.800 59.400 166.200 ;
        RECT 58.200 164.800 58.600 165.200 ;
        RECT 59.000 162.200 59.300 165.800 ;
        RECT 61.400 164.800 61.800 165.200 ;
        RECT 61.400 162.200 61.700 164.800 ;
        RECT 55.800 161.800 56.200 162.200 ;
        RECT 59.000 161.800 59.400 162.200 ;
        RECT 61.400 161.800 61.800 162.200 ;
        RECT 55.000 159.800 55.400 160.200 ;
        RECT 44.600 153.800 45.000 154.200 ;
        RECT 39.800 146.800 40.200 147.200 ;
        RECT 38.200 135.800 38.600 136.200 ;
        RECT 38.200 134.200 38.500 135.800 ;
        RECT 39.000 134.800 39.400 135.200 ;
        RECT 38.200 133.800 38.600 134.200 ;
        RECT 39.000 129.200 39.300 134.800 ;
        RECT 35.000 125.800 35.400 126.200 ;
        RECT 35.800 126.100 36.200 126.200 ;
        RECT 36.600 126.100 37.000 126.200 ;
        RECT 35.800 125.800 37.000 126.100 ;
        RECT 37.400 125.800 37.800 126.200 ;
        RECT 37.400 125.200 37.700 125.800 ;
        RECT 37.400 124.800 37.800 125.200 ;
        RECT 38.200 123.100 38.600 128.900 ;
        RECT 39.000 128.800 39.400 129.200 ;
        RECT 39.800 118.200 40.100 146.800 ;
        RECT 41.400 145.100 41.800 147.900 ;
        RECT 43.000 143.100 43.400 148.900 ;
        RECT 44.600 147.200 44.900 153.800 ;
        RECT 47.000 152.100 47.400 157.900 ;
        RECT 52.600 156.800 53.000 157.200 ;
        RECT 52.600 156.200 52.900 156.800 ;
        RECT 52.600 155.800 53.000 156.200 ;
        RECT 51.800 155.100 52.200 155.200 ;
        RECT 52.600 155.100 53.000 155.200 ;
        RECT 51.800 154.800 53.000 155.100 ;
        RECT 51.800 153.800 52.200 154.200 ;
        RECT 55.000 153.800 55.400 154.200 ;
        RECT 49.400 151.800 49.800 152.200 ;
        RECT 44.600 146.800 45.000 147.200 ;
        RECT 46.200 146.800 46.600 147.200 ;
        RECT 46.200 146.200 46.500 146.800 ;
        RECT 46.200 145.800 46.600 146.200 ;
        RECT 47.800 143.100 48.200 148.900 ;
        RECT 49.400 148.200 49.700 151.800 ;
        RECT 49.400 147.800 49.800 148.200 ;
        RECT 51.800 146.200 52.100 153.800 ;
        RECT 55.000 148.200 55.300 153.800 ;
        RECT 55.800 150.200 56.100 161.800 ;
        RECT 63.000 159.200 63.300 166.800 ;
        RECT 64.600 166.200 64.900 166.800 ;
        RECT 63.800 165.800 64.200 166.200 ;
        RECT 64.600 165.800 65.000 166.200 ;
        RECT 63.000 158.800 63.400 159.200 ;
        RECT 56.600 156.100 57.000 156.200 ;
        RECT 57.400 156.100 57.800 156.200 ;
        RECT 56.600 155.800 57.800 156.100 ;
        RECT 56.600 155.100 57.000 155.200 ;
        RECT 57.400 155.100 57.800 155.200 ;
        RECT 56.600 154.800 57.800 155.100 ;
        RECT 59.800 154.800 60.200 155.200 ;
        RECT 55.800 149.800 56.200 150.200 ;
        RECT 53.400 148.100 53.800 148.200 ;
        RECT 54.200 148.100 54.600 148.200 ;
        RECT 53.400 147.800 54.600 148.100 ;
        RECT 55.000 147.800 55.400 148.200 ;
        RECT 57.400 147.200 57.700 154.800 ;
        RECT 59.800 154.200 60.100 154.800 ;
        RECT 58.200 154.100 58.600 154.200 ;
        RECT 59.000 154.100 59.400 154.200 ;
        RECT 58.200 153.800 59.400 154.100 ;
        RECT 59.800 153.800 60.200 154.200 ;
        RECT 59.800 152.800 60.200 153.200 ;
        RECT 60.600 153.100 61.000 155.900 ;
        RECT 61.400 155.800 61.800 156.200 ;
        RECT 59.800 152.200 60.100 152.800 ;
        RECT 59.800 151.800 60.200 152.200 ;
        RECT 61.400 149.200 61.700 155.800 ;
        RECT 62.200 152.100 62.600 157.900 ;
        RECT 63.000 155.800 63.400 156.200 ;
        RECT 63.000 155.100 63.300 155.800 ;
        RECT 63.000 154.700 63.400 155.100 ;
        RECT 61.400 148.800 61.800 149.200 ;
        RECT 63.000 148.800 63.400 149.200 ;
        RECT 63.000 148.200 63.300 148.800 ;
        RECT 63.000 147.800 63.400 148.200 ;
        RECT 63.800 147.200 64.100 165.800 ;
        RECT 64.600 154.200 64.900 165.800 ;
        RECT 66.200 155.200 66.500 172.800 ;
        RECT 68.600 171.800 69.000 172.200 ;
        RECT 69.400 172.100 69.800 177.900 ;
        RECT 70.200 173.800 70.600 174.200 ;
        RECT 68.600 168.200 68.900 171.800 ;
        RECT 68.600 167.800 69.000 168.200 ;
        RECT 67.000 166.100 67.400 166.200 ;
        RECT 67.800 166.100 68.200 166.200 ;
        RECT 67.000 165.800 68.200 166.100 ;
        RECT 66.200 154.800 66.600 155.200 ;
        RECT 64.600 153.800 65.000 154.200 ;
        RECT 54.200 146.800 54.600 147.200 ;
        RECT 55.800 147.100 56.200 147.200 ;
        RECT 56.600 147.100 57.000 147.200 ;
        RECT 55.800 146.800 57.000 147.100 ;
        RECT 57.400 146.800 57.800 147.200 ;
        RECT 58.200 147.100 58.600 147.200 ;
        RECT 59.000 147.100 59.400 147.200 ;
        RECT 58.200 146.800 59.400 147.100 ;
        RECT 63.800 146.800 64.200 147.200 ;
        RECT 51.800 145.800 52.200 146.200 ;
        RECT 54.200 145.200 54.500 146.800 ;
        RECT 58.200 145.800 58.600 146.200 ;
        RECT 51.800 144.800 52.200 145.200 ;
        RECT 54.200 144.800 54.600 145.200 ;
        RECT 55.800 144.800 56.200 145.200 ;
        RECT 51.800 142.200 52.100 144.800 ;
        RECT 55.800 143.200 56.100 144.800 ;
        RECT 58.200 143.200 58.500 145.800 ;
        RECT 59.000 144.200 59.300 146.800 ;
        RECT 64.600 146.200 64.900 153.800 ;
        RECT 65.400 151.800 65.800 152.200 ;
        RECT 65.400 149.200 65.700 151.800 ;
        RECT 65.400 148.800 65.800 149.200 ;
        RECT 66.200 148.200 66.500 154.800 ;
        RECT 67.000 152.100 67.400 157.900 ;
        RECT 67.000 150.800 67.400 151.200 ;
        RECT 67.000 148.200 67.300 150.800 ;
        RECT 66.200 147.800 66.600 148.200 ;
        RECT 67.000 147.800 67.400 148.200 ;
        RECT 59.800 145.800 60.200 146.200 ;
        RECT 64.600 145.800 65.000 146.200 ;
        RECT 59.800 145.200 60.100 145.800 ;
        RECT 59.800 144.800 60.200 145.200 ;
        RECT 59.000 143.800 59.400 144.200 ;
        RECT 55.800 142.800 56.200 143.200 ;
        RECT 58.200 142.800 58.600 143.200 ;
        RECT 51.800 141.800 52.200 142.200 ;
        RECT 52.600 141.800 53.000 142.200 ;
        RECT 46.200 136.800 46.600 137.200 ;
        RECT 40.600 135.800 41.000 136.200 ;
        RECT 44.600 135.800 45.000 136.200 ;
        RECT 40.600 133.200 40.900 135.800 ;
        RECT 41.400 135.100 41.800 135.200 ;
        RECT 42.200 135.100 42.600 135.200 ;
        RECT 41.400 134.800 42.600 135.100 ;
        RECT 41.400 134.100 41.800 134.200 ;
        RECT 42.200 134.100 42.600 134.200 ;
        RECT 41.400 133.800 42.600 134.100 ;
        RECT 40.600 132.800 41.000 133.200 ;
        RECT 42.200 132.800 42.600 133.200 ;
        RECT 43.800 132.800 44.200 133.200 ;
        RECT 40.600 131.800 41.000 132.200 ;
        RECT 40.600 126.200 40.900 131.800 ;
        RECT 42.200 129.200 42.500 132.800 ;
        RECT 43.000 131.800 43.400 132.200 ;
        RECT 43.000 131.200 43.300 131.800 ;
        RECT 43.000 130.800 43.400 131.200 ;
        RECT 43.800 129.200 44.100 132.800 ;
        RECT 44.600 132.200 44.900 135.800 ;
        RECT 46.200 135.200 46.500 136.800 ;
        RECT 46.200 134.800 46.600 135.200 ;
        RECT 47.000 134.800 47.400 135.200 ;
        RECT 49.400 135.100 49.800 135.200 ;
        RECT 50.200 135.100 50.600 135.200 ;
        RECT 49.400 134.800 50.600 135.100 ;
        RECT 47.000 134.200 47.300 134.800 ;
        RECT 51.800 134.200 52.100 141.800 ;
        RECT 52.600 137.200 52.900 141.800 ;
        RECT 52.600 136.800 53.000 137.200 ;
        RECT 45.400 133.800 45.800 134.200 ;
        RECT 47.000 133.800 47.400 134.200 ;
        RECT 47.800 133.800 48.200 134.200 ;
        RECT 51.800 133.800 52.200 134.200 ;
        RECT 45.400 133.200 45.700 133.800 ;
        RECT 45.400 132.800 45.800 133.200 ;
        RECT 44.600 131.800 45.000 132.200 ;
        RECT 44.600 131.200 44.900 131.800 ;
        RECT 44.600 130.800 45.000 131.200 ;
        RECT 44.600 129.800 45.000 130.200 ;
        RECT 42.200 128.800 42.600 129.200 ;
        RECT 43.000 128.800 43.400 129.200 ;
        RECT 43.800 128.800 44.200 129.200 ;
        RECT 41.400 126.800 41.800 127.200 ;
        RECT 40.600 125.800 41.000 126.200 ;
        RECT 41.400 124.200 41.700 126.800 ;
        RECT 43.000 125.200 43.300 128.800 ;
        RECT 43.800 127.800 44.200 128.200 ;
        RECT 43.800 127.200 44.100 127.800 ;
        RECT 43.800 126.800 44.200 127.200 ;
        RECT 43.000 124.800 43.400 125.200 ;
        RECT 41.400 123.800 41.800 124.200 ;
        RECT 29.400 115.100 29.800 115.200 ;
        RECT 30.200 115.100 30.600 115.200 ;
        RECT 29.400 114.800 30.600 115.100 ;
        RECT 32.600 112.100 33.000 117.900 ;
        RECT 39.800 117.800 40.200 118.200 ;
        RECT 35.800 116.800 36.200 117.200 ;
        RECT 35.800 114.200 36.100 116.800 ;
        RECT 37.400 115.800 37.800 116.200 ;
        RECT 35.800 113.800 36.200 114.200 ;
        RECT 37.400 113.200 37.700 115.800 ;
        RECT 41.400 115.200 41.700 123.800 ;
        RECT 43.000 117.200 43.300 124.800 ;
        RECT 43.800 122.200 44.100 126.800 ;
        RECT 44.600 126.200 44.900 129.800 ;
        RECT 45.400 129.100 45.800 129.200 ;
        RECT 46.200 129.100 46.600 129.200 ;
        RECT 45.400 128.800 46.600 129.100 ;
        RECT 47.000 128.200 47.300 133.800 ;
        RECT 47.800 133.200 48.100 133.800 ;
        RECT 47.800 132.800 48.200 133.200 ;
        RECT 52.600 133.100 53.000 135.900 ;
        RECT 48.600 131.800 49.000 132.200 ;
        RECT 52.600 131.800 53.000 132.200 ;
        RECT 54.200 132.100 54.600 137.900 ;
        RECT 55.800 135.100 56.200 135.200 ;
        RECT 56.600 135.100 57.000 135.200 ;
        RECT 55.800 134.800 57.000 135.100 ;
        RECT 55.000 132.800 55.400 133.200 ;
        RECT 55.800 132.800 56.200 133.200 ;
        RECT 47.000 127.800 47.400 128.200 ;
        RECT 48.600 127.200 48.900 131.800 ;
        RECT 49.400 129.800 49.800 130.200 ;
        RECT 49.400 129.200 49.700 129.800 ;
        RECT 49.400 128.800 49.800 129.200 ;
        RECT 50.200 127.800 50.600 128.200 ;
        RECT 50.200 127.200 50.500 127.800 ;
        RECT 47.000 127.100 47.400 127.200 ;
        RECT 47.800 127.100 48.200 127.200 ;
        RECT 47.000 126.800 48.200 127.100 ;
        RECT 48.600 126.800 49.000 127.200 ;
        RECT 50.200 126.800 50.600 127.200 ;
        RECT 44.600 125.800 45.000 126.200 ;
        RECT 47.800 125.800 48.200 126.200 ;
        RECT 49.400 125.800 49.800 126.200 ;
        RECT 51.000 126.100 51.400 126.200 ;
        RECT 51.800 126.100 52.200 126.200 ;
        RECT 51.000 125.800 52.200 126.100 ;
        RECT 46.200 124.800 46.600 125.200 ;
        RECT 46.200 124.200 46.500 124.800 ;
        RECT 46.200 123.800 46.600 124.200 ;
        RECT 47.800 123.200 48.100 125.800 ;
        RECT 49.400 123.200 49.700 125.800 ;
        RECT 44.600 122.800 45.000 123.200 ;
        RECT 47.800 122.800 48.200 123.200 ;
        RECT 49.400 122.800 49.800 123.200 ;
        RECT 43.800 121.800 44.200 122.200 ;
        RECT 43.000 116.800 43.400 117.200 ;
        RECT 42.200 115.800 42.600 116.200 ;
        RECT 43.800 115.800 44.200 116.200 ;
        RECT 42.200 115.200 42.500 115.800 ;
        RECT 43.800 115.200 44.100 115.800 ;
        RECT 38.200 114.800 38.600 115.200 ;
        RECT 39.800 114.800 40.200 115.200 ;
        RECT 41.400 114.800 41.800 115.200 ;
        RECT 42.200 114.800 42.600 115.200 ;
        RECT 43.800 114.800 44.200 115.200 ;
        RECT 38.200 114.200 38.500 114.800 ;
        RECT 38.200 113.800 38.600 114.200 ;
        RECT 37.400 112.800 37.800 113.200 ;
        RECT 35.000 111.800 35.400 112.200 ;
        RECT 35.000 108.200 35.300 111.800 ;
        RECT 39.800 110.200 40.100 114.800 ;
        RECT 40.600 113.800 41.000 114.200 ;
        RECT 41.400 114.100 41.800 114.200 ;
        RECT 42.200 114.100 42.600 114.200 ;
        RECT 41.400 113.800 42.600 114.100 ;
        RECT 40.600 113.200 40.900 113.800 ;
        RECT 40.600 112.800 41.000 113.200 ;
        RECT 39.800 109.800 40.200 110.200 ;
        RECT 44.600 109.200 44.900 122.800 ;
        RECT 47.000 121.800 47.400 122.200 ;
        RECT 46.200 117.800 46.600 118.200 ;
        RECT 46.200 114.200 46.500 117.800 ;
        RECT 47.000 115.200 47.300 121.800 ;
        RECT 52.600 115.200 52.900 131.800 ;
        RECT 55.000 131.100 55.300 132.800 ;
        RECT 54.200 130.800 55.300 131.100 ;
        RECT 55.800 131.200 56.100 132.800 ;
        RECT 59.000 132.100 59.400 137.900 ;
        RECT 59.800 132.200 60.100 144.800 ;
        RECT 63.800 141.800 64.200 142.200 ;
        RECT 62.200 136.800 62.600 137.200 ;
        RECT 63.800 137.100 64.100 141.800 ;
        RECT 63.800 136.800 64.900 137.100 ;
        RECT 62.200 134.200 62.500 136.800 ;
        RECT 63.800 135.800 64.200 136.200 ;
        RECT 63.800 134.200 64.100 135.800 ;
        RECT 62.200 133.800 62.600 134.200 ;
        RECT 63.800 133.800 64.200 134.200 ;
        RECT 59.800 131.800 60.200 132.200 ;
        RECT 61.400 131.800 61.800 132.200 ;
        RECT 55.800 130.800 56.200 131.200 ;
        RECT 53.400 126.800 53.800 127.200 ;
        RECT 53.400 124.200 53.700 126.800 ;
        RECT 54.200 125.200 54.500 130.800 ;
        RECT 55.000 128.100 55.400 128.200 ;
        RECT 55.800 128.100 56.100 130.800 ;
        RECT 55.000 127.800 56.100 128.100 ;
        RECT 57.400 128.800 57.800 129.200 ;
        RECT 57.400 126.200 57.700 128.800 ;
        RECT 61.400 128.200 61.700 131.800 ;
        RECT 59.000 128.100 59.400 128.200 ;
        RECT 59.800 128.100 60.200 128.200 ;
        RECT 59.000 127.800 60.200 128.100 ;
        RECT 60.600 127.800 61.000 128.200 ;
        RECT 61.400 127.800 61.800 128.200 ;
        RECT 60.600 127.200 60.900 127.800 ;
        RECT 58.200 127.100 58.600 127.200 ;
        RECT 59.000 127.100 59.400 127.200 ;
        RECT 58.200 126.800 59.400 127.100 ;
        RECT 60.600 126.800 61.000 127.200 ;
        RECT 64.600 126.200 64.900 136.800 ;
        RECT 65.400 135.800 65.800 136.200 ;
        RECT 66.200 135.800 66.600 136.200 ;
        RECT 65.400 135.200 65.700 135.800 ;
        RECT 66.200 135.200 66.500 135.800 ;
        RECT 67.000 135.200 67.300 147.800 ;
        RECT 67.800 141.800 68.200 142.200 ;
        RECT 67.800 141.200 68.100 141.800 ;
        RECT 67.800 140.800 68.200 141.200 ;
        RECT 68.600 136.200 68.900 167.800 ;
        RECT 69.400 165.100 69.800 167.900 ;
        RECT 70.200 167.200 70.500 173.800 ;
        RECT 71.000 173.100 71.400 175.900 ;
        RECT 71.000 172.100 71.400 172.200 ;
        RECT 71.800 172.100 72.200 172.200 ;
        RECT 74.200 172.100 74.600 177.900 ;
        RECT 77.400 174.800 77.800 175.200 ;
        RECT 77.400 174.200 77.700 174.800 ;
        RECT 75.000 173.800 75.400 174.200 ;
        RECT 77.400 173.800 77.800 174.200 ;
        RECT 71.000 171.800 72.200 172.100 ;
        RECT 70.200 166.800 70.600 167.200 ;
        RECT 71.000 163.100 71.400 168.900 ;
        RECT 71.800 165.900 72.200 166.300 ;
        RECT 75.000 166.200 75.300 173.800 ;
        RECT 79.000 172.100 79.400 177.900 ;
        RECT 79.800 174.800 80.200 175.200 ;
        RECT 79.800 174.200 80.100 174.800 ;
        RECT 79.800 173.800 80.200 174.200 ;
        RECT 80.600 173.100 81.000 175.900 ;
        RECT 94.200 174.800 94.600 175.200 ;
        RECT 94.200 174.200 94.500 174.800 ;
        RECT 84.600 174.100 85.000 174.200 ;
        RECT 85.400 174.100 85.800 174.200 ;
        RECT 84.600 173.800 85.800 174.100 ;
        RECT 91.000 173.800 91.400 174.200 ;
        RECT 94.200 173.800 94.600 174.200 ;
        RECT 82.200 171.800 82.600 172.200 ;
        RECT 82.200 171.200 82.500 171.800 ;
        RECT 82.200 170.800 82.600 171.200 ;
        RECT 71.000 161.800 71.400 162.200 ;
        RECT 71.000 156.200 71.300 161.800 ;
        RECT 71.000 155.800 71.400 156.200 ;
        RECT 71.000 155.200 71.300 155.800 ;
        RECT 71.800 155.200 72.100 165.900 ;
        RECT 75.000 165.800 75.400 166.200 ;
        RECT 75.800 163.100 76.200 168.900 ;
        RECT 79.000 167.100 79.400 167.200 ;
        RECT 81.400 167.100 81.800 167.200 ;
        RECT 82.200 167.100 82.600 167.200 ;
        RECT 79.000 166.800 80.100 167.100 ;
        RECT 81.400 166.800 82.600 167.100 ;
        RECT 83.800 166.800 84.200 167.200 ;
        RECT 79.000 165.800 79.400 166.200 ;
        RECT 79.000 165.200 79.300 165.800 ;
        RECT 79.000 164.800 79.400 165.200 ;
        RECT 79.800 162.200 80.100 166.800 ;
        RECT 82.200 164.800 82.600 165.200 ;
        RECT 82.200 162.200 82.500 164.800 ;
        RECT 83.800 164.200 84.100 166.800 ;
        RECT 83.800 163.800 84.200 164.200 ;
        RECT 86.200 163.800 86.600 164.200 ;
        RECT 75.800 161.800 76.200 162.200 ;
        RECT 78.200 161.800 78.600 162.200 ;
        RECT 79.800 161.800 80.200 162.200 ;
        RECT 82.200 161.800 82.600 162.200 ;
        RECT 75.000 160.800 75.400 161.200 ;
        RECT 73.400 156.100 73.800 156.200 ;
        RECT 74.200 156.100 74.600 156.200 ;
        RECT 73.400 155.800 74.600 156.100 ;
        RECT 71.000 154.800 71.400 155.200 ;
        RECT 71.800 154.800 72.200 155.200 ;
        RECT 75.000 154.200 75.300 160.800 ;
        RECT 75.800 157.200 76.100 161.800 ;
        RECT 78.200 161.200 78.500 161.800 ;
        RECT 78.200 160.800 78.600 161.200 ;
        RECT 83.800 159.200 84.100 163.800 ;
        RECT 75.800 156.800 76.200 157.200 ;
        RECT 77.400 156.800 77.800 157.200 ;
        RECT 75.800 154.200 76.100 156.800 ;
        RECT 77.400 156.200 77.700 156.800 ;
        RECT 77.400 155.800 77.800 156.200 ;
        RECT 81.400 154.800 81.800 155.200 ;
        RECT 70.200 153.800 70.600 154.200 ;
        RECT 75.000 153.800 75.400 154.200 ;
        RECT 75.800 153.800 76.200 154.200 ;
        RECT 76.600 154.100 77.000 154.200 ;
        RECT 77.400 154.100 77.800 154.200 ;
        RECT 76.600 153.800 77.800 154.100 ;
        RECT 69.400 151.800 69.800 152.200 ;
        RECT 69.400 151.200 69.700 151.800 ;
        RECT 69.400 150.800 69.800 151.200 ;
        RECT 70.200 138.200 70.500 153.800 ;
        RECT 75.000 151.200 75.300 153.800 ;
        RECT 75.000 150.800 75.400 151.200 ;
        RECT 71.800 149.800 72.200 150.200 ;
        RECT 71.800 146.200 72.100 149.800 ;
        RECT 71.800 145.800 72.200 146.200 ;
        RECT 72.600 142.100 73.000 148.900 ;
        RECT 73.400 142.100 73.800 148.900 ;
        RECT 74.200 142.100 74.600 148.900 ;
        RECT 75.000 143.100 75.400 148.900 ;
        RECT 75.800 148.800 76.200 149.200 ;
        RECT 75.800 148.200 76.100 148.800 ;
        RECT 75.800 147.800 76.200 148.200 ;
        RECT 76.600 143.100 77.000 148.900 ;
        RECT 77.400 146.800 77.800 147.200 ;
        RECT 70.200 137.800 70.600 138.200 ;
        RECT 68.600 135.800 69.000 136.200 ;
        RECT 70.200 135.800 70.600 136.200 ;
        RECT 71.000 135.800 71.400 136.200 ;
        RECT 73.400 135.800 73.800 136.200 ;
        RECT 70.200 135.200 70.500 135.800 ;
        RECT 65.400 134.800 65.800 135.200 ;
        RECT 66.200 134.800 66.600 135.200 ;
        RECT 67.000 134.800 67.400 135.200 ;
        RECT 70.200 134.800 70.600 135.200 ;
        RECT 71.000 134.200 71.300 135.800 ;
        RECT 73.400 135.200 73.700 135.800 ;
        RECT 77.400 135.200 77.700 146.800 ;
        RECT 78.200 143.100 78.600 148.900 ;
        RECT 79.000 142.100 79.400 148.900 ;
        RECT 79.800 142.100 80.200 148.900 ;
        RECT 81.400 146.200 81.700 154.800 ;
        RECT 82.200 152.100 82.600 158.900 ;
        RECT 83.000 152.100 83.400 158.900 ;
        RECT 83.800 158.800 84.200 159.200 ;
        RECT 83.800 152.100 84.200 157.900 ;
        RECT 84.600 154.800 85.000 155.200 ;
        RECT 84.600 154.200 84.900 154.800 ;
        RECT 84.600 153.800 85.000 154.200 ;
        RECT 85.400 152.100 85.800 157.900 ;
        RECT 86.200 153.200 86.500 163.800 ;
        RECT 87.000 163.100 87.400 168.900 ;
        RECT 90.200 166.800 90.600 167.200 ;
        RECT 90.200 166.200 90.500 166.800 ;
        RECT 90.200 165.800 90.600 166.200 ;
        RECT 91.000 165.100 91.300 173.800 ;
        RECT 92.600 172.800 93.000 173.200 ;
        RECT 90.200 164.800 91.300 165.100 ;
        RECT 86.200 152.800 86.600 153.200 ;
        RECT 86.200 149.200 86.500 152.800 ;
        RECT 87.000 152.100 87.400 157.900 ;
        RECT 87.800 152.100 88.200 158.900 ;
        RECT 88.600 152.100 89.000 158.900 ;
        RECT 89.400 152.100 89.800 158.900 ;
        RECT 90.200 155.200 90.500 164.800 ;
        RECT 91.800 163.100 92.200 168.900 ;
        RECT 92.600 167.200 92.900 172.800 ;
        RECT 96.600 172.100 97.000 178.900 ;
        RECT 97.400 172.100 97.800 178.900 ;
        RECT 98.200 172.100 98.600 177.900 ;
        RECT 99.000 173.800 99.400 174.200 ;
        RECT 99.000 169.200 99.300 173.800 ;
        RECT 99.800 172.100 100.200 177.900 ;
        RECT 100.600 173.800 101.000 174.200 ;
        RECT 100.600 173.200 100.900 173.800 ;
        RECT 100.600 172.800 101.000 173.200 ;
        RECT 101.400 172.100 101.800 177.900 ;
        RECT 102.200 172.100 102.600 178.900 ;
        RECT 103.000 172.100 103.400 178.900 ;
        RECT 103.800 172.100 104.200 178.900 ;
        RECT 111.800 174.800 112.200 175.200 ;
        RECT 114.200 174.800 114.600 175.200 ;
        RECT 135.000 174.800 135.400 175.200 ;
        RECT 109.400 172.800 109.800 173.200 ;
        RECT 96.600 169.100 97.000 169.200 ;
        RECT 97.400 169.100 97.800 169.200 ;
        RECT 96.600 168.800 97.800 169.100 ;
        RECT 99.000 168.800 99.400 169.200 ;
        RECT 109.400 168.200 109.700 172.800 ;
        RECT 111.800 172.200 112.100 174.800 ;
        RECT 114.200 174.200 114.500 174.800 ;
        RECT 135.000 174.200 135.300 174.800 ;
        RECT 114.200 173.800 114.600 174.200 ;
        RECT 115.000 173.800 115.400 174.200 ;
        RECT 129.400 173.800 129.800 174.200 ;
        RECT 135.000 173.800 135.400 174.200 ;
        RECT 115.000 173.200 115.300 173.800 ;
        RECT 129.400 173.200 129.700 173.800 ;
        RECT 115.000 172.800 115.400 173.200 ;
        RECT 121.400 172.800 121.800 173.200 ;
        RECT 122.200 173.100 122.600 173.200 ;
        RECT 123.000 173.100 123.400 173.200 ;
        RECT 122.200 172.800 123.400 173.100 ;
        RECT 125.400 172.800 125.800 173.200 ;
        RECT 129.400 172.800 129.800 173.200 ;
        RECT 111.800 171.800 112.200 172.200 ;
        RECT 119.000 171.800 119.400 172.200 ;
        RECT 92.600 166.800 93.000 167.200 ;
        RECT 93.400 165.100 93.800 167.900 ;
        RECT 94.900 167.500 95.300 167.900 ;
        RECT 95.800 167.500 97.900 167.800 ;
        RECT 98.200 167.500 98.600 167.900 ;
        RECT 94.200 166.800 94.600 167.200 ;
        RECT 94.200 165.200 94.500 166.800 ;
        RECT 94.200 164.800 94.600 165.200 ;
        RECT 94.900 165.100 95.200 167.500 ;
        RECT 95.800 167.400 96.200 167.500 ;
        RECT 97.500 167.400 97.900 167.500 ;
        RECT 98.300 167.100 98.600 167.500 ;
        RECT 96.200 166.800 98.600 167.100 ;
        RECT 99.000 167.800 99.400 168.200 ;
        RECT 100.600 167.800 101.000 168.200 ;
        RECT 104.600 167.800 105.000 168.200 ;
        RECT 109.400 167.800 109.800 168.200 ;
        RECT 99.000 167.200 99.300 167.800 ;
        RECT 100.600 167.200 100.900 167.800 ;
        RECT 104.600 167.200 104.900 167.800 ;
        RECT 99.000 166.800 99.400 167.200 ;
        RECT 100.600 166.800 101.000 167.200 ;
        RECT 104.600 167.100 105.000 167.200 ;
        RECT 103.800 166.800 105.000 167.100 ;
        RECT 105.400 166.800 105.800 167.200 ;
        RECT 107.000 166.800 107.400 167.200 ;
        RECT 114.200 166.800 114.600 167.200 ;
        RECT 115.800 166.800 116.200 167.200 ;
        RECT 117.400 167.100 117.800 167.200 ;
        RECT 118.200 167.100 118.600 167.200 ;
        RECT 117.400 166.800 118.600 167.100 ;
        RECT 96.200 166.700 96.600 166.800 ;
        RECT 98.300 165.100 98.600 166.800 ;
        RECT 94.900 164.700 95.300 165.100 ;
        RECT 98.200 164.700 98.600 165.100 ;
        RECT 99.000 165.800 99.400 166.200 ;
        RECT 98.200 163.800 98.600 164.200 ;
        RECT 97.400 157.800 97.800 158.200 ;
        RECT 97.400 157.200 97.700 157.800 ;
        RECT 97.400 156.800 97.800 157.200 ;
        RECT 95.800 155.800 96.200 156.200 ;
        RECT 90.200 154.800 90.600 155.200 ;
        RECT 95.800 154.200 96.100 155.800 ;
        RECT 98.200 154.200 98.500 163.800 ;
        RECT 99.000 155.200 99.300 165.800 ;
        RECT 103.000 161.800 103.400 162.200 ;
        RECT 103.000 161.200 103.300 161.800 ;
        RECT 103.000 160.800 103.400 161.200 ;
        RECT 103.800 159.200 104.100 166.800 ;
        RECT 103.800 158.800 104.200 159.200 ;
        RECT 99.000 154.800 99.400 155.200 ;
        RECT 95.800 153.800 96.200 154.200 ;
        RECT 98.200 153.800 98.600 154.200 ;
        RECT 100.600 153.800 101.000 154.200 ;
        RECT 104.600 153.800 105.000 154.200 ;
        RECT 100.600 153.200 100.900 153.800 ;
        RECT 104.600 153.200 104.900 153.800 ;
        RECT 100.600 152.800 101.000 153.200 ;
        RECT 104.600 152.800 105.000 153.200 ;
        RECT 99.800 151.800 100.200 152.200 ;
        RECT 86.200 148.800 86.600 149.200 ;
        RECT 83.800 148.100 84.200 148.200 ;
        RECT 84.600 148.100 85.000 148.200 ;
        RECT 83.800 147.800 85.000 148.100 ;
        RECT 86.200 146.800 86.600 147.200 ;
        RECT 88.600 147.100 89.000 147.200 ;
        RECT 89.400 147.100 89.800 147.200 ;
        RECT 88.600 146.800 89.800 147.100 ;
        RECT 81.400 145.800 81.800 146.200 ;
        RECT 85.400 141.800 85.800 142.200 ;
        RECT 78.200 139.800 78.600 140.200 ;
        RECT 80.600 139.800 81.000 140.200 ;
        RECT 78.200 136.200 78.500 139.800 ;
        RECT 78.200 135.800 78.600 136.200 ;
        RECT 80.600 135.200 80.900 139.800 ;
        RECT 73.400 134.800 73.800 135.200 ;
        RECT 74.200 134.800 74.600 135.200 ;
        RECT 77.400 134.800 77.800 135.200 ;
        RECT 79.000 135.100 79.400 135.200 ;
        RECT 79.800 135.100 80.200 135.200 ;
        RECT 79.000 134.800 80.200 135.100 ;
        RECT 80.600 134.800 81.000 135.200 ;
        RECT 74.200 134.200 74.500 134.800 ;
        RECT 66.200 134.100 66.600 134.200 ;
        RECT 67.000 134.100 67.400 134.200 ;
        RECT 66.200 133.800 67.400 134.100 ;
        RECT 67.800 133.800 68.200 134.200 ;
        RECT 69.400 133.800 69.800 134.200 ;
        RECT 71.000 133.800 71.400 134.200 ;
        RECT 72.600 133.800 73.000 134.200 ;
        RECT 74.200 133.800 74.600 134.200 ;
        RECT 76.600 133.800 77.000 134.200 ;
        RECT 81.400 133.800 81.800 134.200 ;
        RECT 67.800 132.200 68.100 133.800 ;
        RECT 67.800 131.800 68.200 132.200 ;
        RECT 67.800 127.800 68.200 128.200 ;
        RECT 67.800 127.200 68.100 127.800 ;
        RECT 69.400 127.200 69.700 133.800 ;
        RECT 70.200 131.800 70.600 132.200 ;
        RECT 71.800 131.800 72.200 132.200 ;
        RECT 70.200 129.200 70.500 131.800 ;
        RECT 70.200 128.800 70.600 129.200 ;
        RECT 65.400 126.800 65.800 127.200 ;
        RECT 66.200 127.100 66.600 127.200 ;
        RECT 67.000 127.100 67.400 127.200 ;
        RECT 66.200 126.800 67.400 127.100 ;
        RECT 67.800 126.800 68.200 127.200 ;
        RECT 69.400 126.800 69.800 127.200 ;
        RECT 70.200 126.800 70.600 127.200 ;
        RECT 57.400 125.800 57.800 126.200 ;
        RECT 63.800 125.800 64.200 126.200 ;
        RECT 64.600 125.800 65.000 126.200 ;
        RECT 54.200 124.800 54.600 125.200 ;
        RECT 55.800 124.800 56.200 125.200 ;
        RECT 57.400 125.100 57.800 125.200 ;
        RECT 59.000 125.100 59.400 125.200 ;
        RECT 57.400 124.800 59.400 125.100 ;
        RECT 63.000 124.800 63.400 125.200 ;
        RECT 55.800 124.200 56.100 124.800 ;
        RECT 53.400 123.800 53.800 124.200 ;
        RECT 55.800 123.800 56.200 124.200 ;
        RECT 63.000 123.200 63.300 124.800 ;
        RECT 55.000 122.800 55.400 123.200 ;
        RECT 63.000 122.800 63.400 123.200 ;
        RECT 55.000 122.200 55.300 122.800 ;
        RECT 55.000 121.800 55.400 122.200 ;
        RECT 62.200 121.800 62.600 122.200 ;
        RECT 61.400 118.800 61.800 119.200 ;
        RECT 58.200 117.800 58.600 118.200 ;
        RECT 53.400 115.800 53.800 116.200 ;
        RECT 55.800 115.800 56.200 116.200 ;
        RECT 53.400 115.200 53.700 115.800 ;
        RECT 47.000 114.800 47.400 115.200 ;
        RECT 51.000 114.800 51.400 115.200 ;
        RECT 52.600 114.800 53.000 115.200 ;
        RECT 53.400 114.800 53.800 115.200 ;
        RECT 47.000 114.200 47.300 114.800 ;
        RECT 46.200 113.800 46.600 114.200 ;
        RECT 47.000 113.800 47.400 114.200 ;
        RECT 47.800 114.100 48.200 114.200 ;
        RECT 48.600 114.100 49.000 114.200 ;
        RECT 47.800 113.800 49.000 114.100 ;
        RECT 45.400 111.800 45.800 112.200 ;
        RECT 45.400 111.200 45.700 111.800 ;
        RECT 45.400 110.800 45.800 111.200 ;
        RECT 47.000 110.200 47.300 113.800 ;
        RECT 47.800 113.200 48.100 113.800 ;
        RECT 47.800 112.800 48.200 113.200 ;
        RECT 47.000 109.800 47.400 110.200 ;
        RECT 35.800 108.800 36.200 109.200 ;
        RECT 44.600 108.800 45.000 109.200 ;
        RECT 31.000 108.100 31.400 108.200 ;
        RECT 31.800 108.100 32.200 108.200 ;
        RECT 31.000 107.800 32.200 108.100 ;
        RECT 35.000 107.800 35.400 108.200 ;
        RECT 29.400 107.100 29.800 107.200 ;
        RECT 30.200 107.100 30.600 107.200 ;
        RECT 29.400 106.800 30.600 107.100 ;
        RECT 34.200 107.100 34.600 107.200 ;
        RECT 35.000 107.100 35.400 107.200 ;
        RECT 34.200 106.800 35.400 107.100 ;
        RECT 26.200 106.100 26.600 106.200 ;
        RECT 27.000 106.100 27.400 106.200 ;
        RECT 26.200 105.800 27.400 106.100 ;
        RECT 28.600 105.800 29.000 106.200 ;
        RECT 31.800 106.100 32.200 106.200 ;
        RECT 32.600 106.100 33.000 106.200 ;
        RECT 31.800 105.800 33.000 106.100 ;
        RECT 33.400 105.800 33.800 106.200 ;
        RECT 35.800 106.100 36.100 108.800 ;
        RECT 47.000 108.200 47.300 109.800 ;
        RECT 39.800 108.100 40.200 108.200 ;
        RECT 40.600 108.100 41.000 108.200 ;
        RECT 39.800 107.800 41.000 108.100 ;
        RECT 43.800 107.800 44.200 108.200 ;
        RECT 45.400 108.100 45.800 108.200 ;
        RECT 46.200 108.100 46.600 108.200 ;
        RECT 45.400 107.800 46.600 108.100 ;
        RECT 47.000 107.800 47.400 108.200 ;
        RECT 43.800 107.200 44.100 107.800 ;
        RECT 51.000 107.200 51.300 114.800 ;
        RECT 55.800 114.200 56.100 115.800 ;
        RECT 58.200 114.200 58.500 117.800 ;
        RECT 61.400 115.200 61.700 118.800 ;
        RECT 62.200 115.200 62.500 121.800 ;
        RECT 63.800 119.200 64.100 125.800 ;
        RECT 65.400 124.200 65.700 126.800 ;
        RECT 70.200 126.200 70.500 126.800 ;
        RECT 66.200 126.100 66.600 126.200 ;
        RECT 67.000 126.100 67.400 126.200 ;
        RECT 66.200 125.800 67.400 126.100 ;
        RECT 70.200 125.800 70.600 126.200 ;
        RECT 71.000 125.800 71.400 126.200 ;
        RECT 71.000 125.200 71.300 125.800 ;
        RECT 71.800 125.200 72.100 131.800 ;
        RECT 72.600 129.200 72.900 133.800 ;
        RECT 72.600 128.800 73.000 129.200 ;
        RECT 67.800 124.800 68.200 125.200 ;
        RECT 68.600 124.800 69.000 125.200 ;
        RECT 71.000 124.800 71.400 125.200 ;
        RECT 71.800 124.800 72.200 125.200 ;
        RECT 65.400 123.800 65.800 124.200 ;
        RECT 63.800 118.800 64.200 119.200 ;
        RECT 63.800 118.100 64.200 118.200 ;
        RECT 64.600 118.100 65.000 118.200 ;
        RECT 63.800 117.800 65.000 118.100 ;
        RECT 63.800 116.100 64.200 116.200 ;
        RECT 63.800 115.800 64.900 116.100 ;
        RECT 61.400 114.800 61.800 115.200 ;
        RECT 62.200 114.800 62.600 115.200 ;
        RECT 51.800 114.100 52.200 114.200 ;
        RECT 52.600 114.100 53.000 114.200 ;
        RECT 51.800 113.800 53.000 114.100 ;
        RECT 55.800 113.800 56.200 114.200 ;
        RECT 58.200 113.800 58.600 114.200 ;
        RECT 59.800 114.100 60.200 114.200 ;
        RECT 60.600 114.100 61.000 114.200 ;
        RECT 59.800 113.800 61.000 114.100 ;
        RECT 61.400 113.800 61.800 114.200 ;
        RECT 63.000 114.100 63.400 114.200 ;
        RECT 63.800 114.100 64.200 114.200 ;
        RECT 63.000 113.800 64.200 114.100 ;
        RECT 61.400 113.200 61.700 113.800 ;
        RECT 52.600 112.800 53.000 113.200 ;
        RECT 58.200 112.800 58.600 113.200 ;
        RECT 61.400 112.800 61.800 113.200 ;
        RECT 63.800 112.800 64.200 113.200 ;
        RECT 52.600 109.200 52.900 112.800 ;
        RECT 55.000 111.800 55.400 112.200 ;
        RECT 55.000 111.200 55.300 111.800 ;
        RECT 55.000 110.800 55.400 111.200 ;
        RECT 58.200 110.200 58.500 112.800 ;
        RECT 59.000 111.800 59.400 112.200 ;
        RECT 55.000 109.800 55.400 110.200 ;
        RECT 58.200 109.800 58.600 110.200 ;
        RECT 55.000 109.200 55.300 109.800 ;
        RECT 52.600 108.800 53.000 109.200 ;
        RECT 55.000 108.800 55.400 109.200 ;
        RECT 57.400 109.100 57.800 109.200 ;
        RECT 58.200 109.100 58.600 109.200 ;
        RECT 57.400 108.800 58.600 109.100 ;
        RECT 36.600 107.100 37.000 107.200 ;
        RECT 37.400 107.100 37.800 107.200 ;
        RECT 36.600 106.800 37.800 107.100 ;
        RECT 41.400 107.100 41.800 107.200 ;
        RECT 42.200 107.100 42.600 107.200 ;
        RECT 41.400 106.800 42.600 107.100 ;
        RECT 43.800 106.800 44.200 107.200 ;
        RECT 45.400 107.100 45.800 107.200 ;
        RECT 46.200 107.100 46.600 107.200 ;
        RECT 45.400 106.800 46.600 107.100 ;
        RECT 51.000 106.800 51.400 107.200 ;
        RECT 57.400 106.800 57.800 107.200 ;
        RECT 57.400 106.200 57.700 106.800 ;
        RECT 36.600 106.100 37.000 106.200 ;
        RECT 35.800 105.800 37.000 106.100 ;
        RECT 38.200 105.800 38.600 106.200 ;
        RECT 42.200 105.800 42.600 106.200 ;
        RECT 43.000 105.800 43.400 106.200 ;
        RECT 51.000 106.100 51.400 106.200 ;
        RECT 51.800 106.100 52.200 106.200 ;
        RECT 51.000 105.800 52.200 106.100 ;
        RECT 52.600 105.800 53.000 106.200 ;
        RECT 56.600 105.800 57.000 106.200 ;
        RECT 57.400 105.800 57.800 106.200 ;
        RECT 58.200 105.800 58.600 106.200 ;
        RECT 59.000 106.100 59.300 111.800 ;
        RECT 60.600 106.800 61.000 107.200 ;
        RECT 61.400 106.800 61.800 107.200 ;
        RECT 59.800 106.100 60.200 106.200 ;
        RECT 59.000 105.800 60.200 106.100 ;
        RECT 26.200 105.100 26.600 105.200 ;
        RECT 25.400 104.800 26.600 105.100 ;
        RECT 25.400 99.200 25.700 104.800 ;
        RECT 33.400 104.200 33.700 105.800 ;
        RECT 27.000 103.800 27.400 104.200 ;
        RECT 33.400 103.800 33.800 104.200 ;
        RECT 27.000 99.200 27.300 103.800 ;
        RECT 37.400 102.800 37.800 103.200 ;
        RECT 35.800 101.800 36.200 102.200 ;
        RECT 25.400 98.800 25.800 99.200 ;
        RECT 27.000 98.800 27.400 99.200 ;
        RECT 27.800 98.800 28.200 99.200 ;
        RECT 27.800 95.200 28.100 98.800 ;
        RECT 30.200 97.800 30.600 98.200 ;
        RECT 30.200 97.200 30.500 97.800 ;
        RECT 30.200 96.800 30.600 97.200 ;
        RECT 27.800 94.800 28.200 95.200 ;
        RECT 31.000 94.800 31.400 95.200 ;
        RECT 31.800 94.800 32.200 95.200 ;
        RECT 33.400 95.100 33.800 95.200 ;
        RECT 34.200 95.100 34.600 95.200 ;
        RECT 33.400 94.800 34.600 95.100 ;
        RECT 35.000 95.100 35.400 95.200 ;
        RECT 35.800 95.100 36.100 101.800 ;
        RECT 36.600 96.800 37.000 97.200 ;
        RECT 36.600 96.200 36.900 96.800 ;
        RECT 36.600 95.800 37.000 96.200 ;
        RECT 35.000 94.800 36.100 95.100 ;
        RECT 37.400 95.200 37.700 102.800 ;
        RECT 38.200 99.200 38.500 105.800 ;
        RECT 42.200 105.200 42.500 105.800 ;
        RECT 43.000 105.200 43.300 105.800 ;
        RECT 42.200 104.800 42.600 105.200 ;
        RECT 43.000 104.800 43.400 105.200 ;
        RECT 39.800 103.800 40.200 104.200 ;
        RECT 38.200 98.800 38.600 99.200 ;
        RECT 39.800 96.200 40.100 103.800 ;
        RECT 47.800 99.100 48.200 99.200 ;
        RECT 48.600 99.100 49.000 99.200 ;
        RECT 47.800 98.800 49.000 99.100 ;
        RECT 47.800 97.800 48.200 98.200 ;
        RECT 39.800 95.800 40.200 96.200 ;
        RECT 41.400 95.800 41.800 96.200 ;
        RECT 43.800 95.800 44.200 96.200 ;
        RECT 45.400 95.800 45.800 96.200 ;
        RECT 37.400 94.800 37.800 95.200 ;
        RECT 23.800 94.100 24.200 94.200 ;
        RECT 23.000 93.800 24.200 94.100 ;
        RECT 27.800 93.800 28.200 94.200 ;
        RECT 23.000 88.200 23.300 93.800 ;
        RECT 25.400 92.800 25.800 93.200 ;
        RECT 26.200 93.100 26.600 93.200 ;
        RECT 27.000 93.100 27.400 93.200 ;
        RECT 26.200 92.800 27.400 93.100 ;
        RECT 25.400 89.200 25.700 92.800 ;
        RECT 27.800 91.200 28.100 93.800 ;
        RECT 28.600 92.800 29.000 93.200 ;
        RECT 30.200 92.800 30.600 93.200 ;
        RECT 27.800 90.800 28.200 91.200 ;
        RECT 25.400 88.800 25.800 89.200 ;
        RECT 23.000 87.800 23.400 88.200 ;
        RECT 23.000 86.200 23.300 87.800 ;
        RECT 23.800 86.800 24.200 87.200 ;
        RECT 22.200 85.800 22.600 86.200 ;
        RECT 23.000 85.800 23.400 86.200 ;
        RECT 22.200 79.200 22.500 85.800 ;
        RECT 23.800 80.200 24.100 86.800 ;
        RECT 24.600 85.100 25.000 87.900 ;
        RECT 25.400 87.800 25.800 88.200 ;
        RECT 25.400 87.200 25.700 87.800 ;
        RECT 25.400 86.800 25.800 87.200 ;
        RECT 26.200 83.100 26.600 88.900 ;
        RECT 27.800 87.800 28.200 88.200 ;
        RECT 27.800 86.200 28.100 87.800 ;
        RECT 27.800 85.800 28.200 86.200 ;
        RECT 23.800 79.800 24.200 80.200 ;
        RECT 22.200 78.800 22.600 79.200 ;
        RECT 27.000 79.100 27.400 79.200 ;
        RECT 27.800 79.100 28.200 79.200 ;
        RECT 27.000 78.800 28.200 79.100 ;
        RECT 20.600 72.100 21.000 77.900 ;
        RECT 21.400 75.800 21.800 76.200 ;
        RECT 21.400 75.100 21.700 75.800 ;
        RECT 21.400 74.700 21.800 75.100 ;
        RECT 24.600 73.800 25.000 74.200 ;
        RECT 24.600 73.200 24.900 73.800 ;
        RECT 21.400 72.800 21.800 73.200 ;
        RECT 24.600 72.800 25.000 73.200 ;
        RECT 21.400 67.200 21.700 72.800 ;
        RECT 25.400 72.100 25.800 77.900 ;
        RECT 28.600 74.200 28.900 92.800 ;
        RECT 29.400 90.800 29.800 91.200 ;
        RECT 29.400 87.200 29.700 90.800 ;
        RECT 30.200 90.200 30.500 92.800 ;
        RECT 31.000 90.200 31.300 94.800 ;
        RECT 31.800 94.200 32.100 94.800 ;
        RECT 31.800 93.800 32.200 94.200 ;
        RECT 33.400 93.800 33.800 94.200 ;
        RECT 34.200 93.800 34.600 94.200 ;
        RECT 35.800 93.800 36.200 94.200 ;
        RECT 37.400 93.800 37.800 94.200 ;
        RECT 33.400 93.200 33.700 93.800 ;
        RECT 33.400 92.800 33.800 93.200 ;
        RECT 34.200 90.200 34.500 93.800 ;
        RECT 35.800 93.200 36.100 93.800 ;
        RECT 35.800 92.800 36.200 93.200 ;
        RECT 37.400 90.200 37.700 93.800 ;
        RECT 39.800 93.200 40.100 95.800 ;
        RECT 41.400 95.200 41.700 95.800 ;
        RECT 41.400 94.800 41.800 95.200 ;
        RECT 43.000 94.800 43.400 95.200 ;
        RECT 42.200 94.100 42.600 94.200 ;
        RECT 41.400 93.800 42.600 94.100 ;
        RECT 39.800 92.800 40.200 93.200 ;
        RECT 30.200 89.800 30.600 90.200 ;
        RECT 31.000 89.800 31.400 90.200 ;
        RECT 34.200 89.800 34.600 90.200 ;
        RECT 37.400 89.800 37.800 90.200 ;
        RECT 29.400 86.800 29.800 87.200 ;
        RECT 31.000 83.100 31.400 88.900 ;
        RECT 37.400 88.800 37.800 89.200 ;
        RECT 37.400 88.200 37.700 88.800 ;
        RECT 37.400 87.800 37.800 88.200 ;
        RECT 34.200 86.800 34.600 87.200 ;
        RECT 35.800 86.800 36.200 87.200 ;
        RECT 38.200 87.100 38.600 87.200 ;
        RECT 39.000 87.100 39.400 87.200 ;
        RECT 38.200 86.800 39.400 87.100 ;
        RECT 40.600 86.800 41.000 87.200 ;
        RECT 34.200 86.200 34.500 86.800 ;
        RECT 35.800 86.200 36.100 86.800 ;
        RECT 34.200 85.800 34.600 86.200 ;
        RECT 35.800 85.800 36.200 86.200 ;
        RECT 31.000 79.800 31.400 80.200 ;
        RECT 31.000 79.200 31.300 79.800 ;
        RECT 31.000 78.800 31.400 79.200 ;
        RECT 30.200 76.800 30.600 77.200 ;
        RECT 30.200 76.200 30.500 76.800 ;
        RECT 30.200 75.800 30.600 76.200 ;
        RECT 28.600 73.800 29.000 74.200 ;
        RECT 28.600 70.200 28.900 73.800 ;
        RECT 29.400 71.800 29.800 72.200 ;
        RECT 24.600 69.800 25.000 70.200 ;
        RECT 28.600 69.800 29.000 70.200 ;
        RECT 24.600 69.200 24.900 69.800 ;
        RECT 21.400 66.800 21.800 67.200 ;
        RECT 22.200 63.100 22.600 68.900 ;
        RECT 24.600 68.800 25.000 69.200 ;
        RECT 29.400 68.200 29.700 71.800 ;
        RECT 27.000 67.800 27.400 68.200 ;
        RECT 27.800 67.800 28.200 68.200 ;
        RECT 29.400 67.800 29.800 68.200 ;
        RECT 27.000 67.200 27.300 67.800 ;
        RECT 25.400 67.100 25.800 67.200 ;
        RECT 26.200 67.100 26.600 67.200 ;
        RECT 25.400 66.800 26.600 67.100 ;
        RECT 27.000 66.800 27.400 67.200 ;
        RECT 25.400 66.100 25.800 66.200 ;
        RECT 26.200 66.100 26.600 66.200 ;
        RECT 25.400 65.800 26.600 66.100 ;
        RECT 27.800 65.200 28.100 67.800 ;
        RECT 30.200 67.200 30.500 75.800 ;
        RECT 31.800 72.800 32.200 73.200 ;
        RECT 32.600 73.100 33.000 75.900 ;
        RECT 33.400 74.800 33.800 75.200 ;
        RECT 33.400 74.200 33.700 74.800 ;
        RECT 33.400 73.800 33.800 74.200 ;
        RECT 31.800 72.200 32.100 72.800 ;
        RECT 31.800 71.800 32.200 72.200 ;
        RECT 34.200 72.100 34.600 77.900 ;
        RECT 35.800 75.100 36.200 75.200 ;
        RECT 36.600 75.100 37.000 75.200 ;
        RECT 35.800 74.800 37.000 75.100 ;
        RECT 36.600 73.800 37.000 74.200 ;
        RECT 35.000 72.800 35.400 73.200 ;
        RECT 33.400 67.800 33.800 68.200 ;
        RECT 33.400 67.200 33.700 67.800 ;
        RECT 28.600 66.800 29.000 67.200 ;
        RECT 30.200 66.800 30.600 67.200 ;
        RECT 33.400 66.800 33.800 67.200 ;
        RECT 28.600 65.200 28.900 66.800 ;
        RECT 29.400 66.100 29.800 66.200 ;
        RECT 30.200 66.100 30.600 66.200 ;
        RECT 29.400 65.800 30.600 66.100 ;
        RECT 31.800 66.100 32.200 66.200 ;
        RECT 32.600 66.100 33.000 66.200 ;
        RECT 31.800 65.800 33.000 66.100 ;
        RECT 27.800 64.800 28.200 65.200 ;
        RECT 28.600 64.800 29.000 65.200 ;
        RECT 24.600 57.800 25.000 58.200 ;
        RECT 20.600 57.100 21.000 57.200 ;
        RECT 21.400 57.100 21.800 57.200 ;
        RECT 20.600 56.800 21.800 57.100 ;
        RECT 19.800 55.800 20.200 56.200 ;
        RECT 22.200 56.100 22.600 56.200 ;
        RECT 23.000 56.100 23.400 56.200 ;
        RECT 22.200 55.800 23.400 56.100 ;
        RECT 19.800 55.200 20.100 55.800 ;
        RECT 24.600 55.200 24.900 57.800 ;
        RECT 19.000 54.800 19.400 55.200 ;
        RECT 19.800 54.800 20.200 55.200 ;
        RECT 24.600 54.800 25.000 55.200 ;
        RECT 24.600 54.200 24.900 54.800 ;
        RECT 19.800 53.800 20.200 54.200 ;
        RECT 24.600 53.800 25.000 54.200 ;
        RECT 19.000 46.800 19.400 47.200 ;
        RECT 16.600 46.100 17.000 46.200 ;
        RECT 17.400 46.100 17.800 46.200 ;
        RECT 16.600 45.800 17.800 46.100 ;
        RECT 18.200 45.800 18.600 46.200 ;
        RECT 18.200 45.200 18.500 45.800 ;
        RECT 18.200 44.800 18.600 45.200 ;
        RECT 19.000 44.200 19.300 46.800 ;
        RECT 19.000 43.800 19.400 44.200 ;
        RECT 19.800 37.200 20.100 53.800 ;
        RECT 25.400 53.100 25.800 55.900 ;
        RECT 27.000 52.100 27.400 57.900 ;
        RECT 27.800 52.800 28.200 53.200 ;
        RECT 23.800 48.800 24.200 49.200 ;
        RECT 23.800 47.200 24.100 48.800 ;
        RECT 22.200 46.800 22.600 47.200 ;
        RECT 23.800 46.800 24.200 47.200 ;
        RECT 22.200 46.200 22.500 46.800 ;
        RECT 22.200 45.800 22.600 46.200 ;
        RECT 22.200 45.100 22.600 45.200 ;
        RECT 23.000 45.100 23.400 45.200 ;
        RECT 24.600 45.100 25.000 47.900 ;
        RECT 25.400 46.800 25.800 47.200 ;
        RECT 22.200 44.800 23.400 45.100 ;
        RECT 22.200 43.800 22.600 44.200 ;
        RECT 15.800 36.800 16.200 37.200 ;
        RECT 19.800 36.800 20.200 37.200 ;
        RECT 15.800 35.800 16.200 36.200 ;
        RECT 18.200 35.800 18.600 36.200 ;
        RECT 15.800 35.200 16.100 35.800 ;
        RECT 18.200 35.200 18.500 35.800 ;
        RECT 22.200 35.200 22.500 43.800 ;
        RECT 12.600 35.100 13.000 35.200 ;
        RECT 11.800 34.800 13.000 35.100 ;
        RECT 14.200 35.100 14.600 35.200 ;
        RECT 15.000 35.100 15.400 35.200 ;
        RECT 14.200 34.800 15.400 35.100 ;
        RECT 15.800 34.800 16.200 35.200 ;
        RECT 18.200 34.800 18.600 35.200 ;
        RECT 19.000 34.800 19.400 35.200 ;
        RECT 22.200 34.800 22.600 35.200 ;
        RECT 10.200 32.800 10.600 33.200 ;
        RECT 6.200 26.800 6.600 27.200 ;
        RECT 6.200 26.200 6.500 26.800 ;
        RECT 7.000 26.300 7.300 31.800 ;
        RECT 10.200 29.200 10.500 32.800 ;
        RECT 6.200 25.800 6.600 26.200 ;
        RECT 7.000 25.900 7.400 26.300 ;
        RECT 7.000 25.800 7.300 25.900 ;
        RECT 0.600 13.100 1.000 15.900 ;
        RECT 2.200 12.100 2.600 17.900 ;
        RECT 6.200 15.200 6.500 25.800 ;
        RECT 7.800 23.100 8.200 28.900 ;
        RECT 10.200 28.800 10.600 29.200 ;
        RECT 9.400 25.100 9.800 27.900 ;
        RECT 5.400 14.800 5.800 15.200 ;
        RECT 6.200 14.800 6.600 15.200 ;
        RECT 5.400 13.200 5.700 14.800 ;
        RECT 5.400 12.800 5.800 13.200 ;
        RECT 6.200 9.200 6.500 14.800 ;
        RECT 7.000 12.100 7.400 17.900 ;
        RECT 11.800 16.200 12.100 34.800 ;
        RECT 19.000 34.200 19.300 34.800 ;
        RECT 16.600 34.100 17.000 34.200 ;
        RECT 17.400 34.100 17.800 34.200 ;
        RECT 16.600 33.800 17.800 34.100 ;
        RECT 19.000 33.800 19.400 34.200 ;
        RECT 15.800 33.100 16.200 33.200 ;
        RECT 16.600 33.100 17.000 33.200 ;
        RECT 15.800 32.800 17.000 33.100 ;
        RECT 12.600 32.100 13.000 32.200 ;
        RECT 13.400 32.100 13.800 32.200 ;
        RECT 12.600 31.800 13.800 32.100 ;
        RECT 16.600 31.800 17.000 32.200 ;
        RECT 19.800 32.100 20.200 32.200 ;
        RECT 20.600 32.100 21.000 32.200 ;
        RECT 19.800 31.800 21.000 32.100 ;
        RECT 12.600 23.100 13.000 28.900 ;
        RECT 13.400 26.800 13.800 27.200 ;
        RECT 13.400 26.200 13.700 26.800 ;
        RECT 16.600 26.300 16.900 31.800 ;
        RECT 13.400 25.800 13.800 26.200 ;
        RECT 16.600 25.900 17.000 26.300 ;
        RECT 16.600 25.800 16.900 25.900 ;
        RECT 15.000 22.800 15.400 23.200 ;
        RECT 17.400 23.100 17.800 28.900 ;
        RECT 19.000 25.100 19.400 27.900 ;
        RECT 19.800 25.100 20.200 27.900 ;
        RECT 20.600 26.800 21.000 27.200 ;
        RECT 10.200 15.800 10.600 16.200 ;
        RECT 11.800 15.800 12.200 16.200 ;
        RECT 10.200 15.200 10.500 15.800 ;
        RECT 10.200 14.800 10.600 15.200 ;
        RECT 11.000 14.800 11.400 15.200 ;
        RECT 13.400 15.100 13.800 15.200 ;
        RECT 14.200 15.100 14.600 15.200 ;
        RECT 13.400 14.800 14.600 15.100 ;
        RECT 11.000 14.200 11.300 14.800 ;
        RECT 15.000 14.200 15.300 22.800 ;
        RECT 9.400 14.100 9.800 14.200 ;
        RECT 10.200 14.100 10.600 14.200 ;
        RECT 9.400 13.800 10.600 14.100 ;
        RECT 11.000 13.800 11.400 14.200 ;
        RECT 15.000 13.800 15.400 14.200 ;
        RECT 15.000 13.200 15.300 13.800 ;
        RECT 11.000 13.100 11.400 13.200 ;
        RECT 11.800 13.100 12.200 13.200 ;
        RECT 11.000 12.800 12.200 13.100 ;
        RECT 15.000 12.800 15.400 13.200 ;
        RECT 15.800 13.100 16.200 15.900 ;
        RECT 17.400 12.100 17.800 17.900 ;
        RECT 20.600 15.200 20.900 26.800 ;
        RECT 21.400 23.100 21.800 28.900 ;
        RECT 22.200 26.200 22.500 34.800 ;
        RECT 23.000 33.100 23.400 35.900 ;
        RECT 24.600 32.100 25.000 37.900 ;
        RECT 25.400 33.200 25.700 46.800 ;
        RECT 26.200 43.100 26.600 48.900 ;
        RECT 27.800 47.200 28.100 52.800 ;
        RECT 27.800 46.800 28.200 47.200 ;
        RECT 27.000 46.200 27.400 46.300 ;
        RECT 27.800 46.200 28.200 46.300 ;
        RECT 27.000 45.900 28.200 46.200 ;
        RECT 28.600 36.200 28.900 64.800 ;
        RECT 30.200 62.200 30.500 65.800 ;
        RECT 31.000 64.800 31.400 65.200 ;
        RECT 31.800 65.100 32.200 65.200 ;
        RECT 32.600 65.100 33.000 65.200 ;
        RECT 34.200 65.100 34.600 67.900 ;
        RECT 31.800 64.800 33.000 65.100 ;
        RECT 31.000 64.200 31.300 64.800 ;
        RECT 31.000 63.800 31.400 64.200 ;
        RECT 32.600 64.100 33.000 64.200 ;
        RECT 33.400 64.100 33.800 64.200 ;
        RECT 32.600 63.800 33.800 64.100 ;
        RECT 30.200 61.800 30.600 62.200 ;
        RECT 29.400 55.100 29.800 55.200 ;
        RECT 30.200 55.100 30.600 55.200 ;
        RECT 29.400 54.800 30.600 55.100 ;
        RECT 31.800 52.100 32.200 57.900 ;
        RECT 35.000 57.200 35.300 72.800 ;
        RECT 35.800 63.100 36.200 68.900 ;
        RECT 36.600 68.200 36.900 73.800 ;
        RECT 36.600 67.800 37.000 68.200 ;
        RECT 36.600 66.100 37.000 66.300 ;
        RECT 37.400 66.100 37.800 66.200 ;
        RECT 36.600 65.800 37.800 66.100 ;
        RECT 38.200 59.200 38.500 86.800 ;
        RECT 40.600 86.200 40.900 86.800 ;
        RECT 39.000 85.800 39.400 86.200 ;
        RECT 39.800 85.800 40.200 86.200 ;
        RECT 40.600 85.800 41.000 86.200 ;
        RECT 39.000 84.200 39.300 85.800 ;
        RECT 39.800 85.200 40.100 85.800 ;
        RECT 39.800 84.800 40.200 85.200 ;
        RECT 39.000 83.800 39.400 84.200 ;
        RECT 41.400 82.200 41.700 93.800 ;
        RECT 42.200 92.800 42.600 93.200 ;
        RECT 42.200 92.200 42.500 92.800 ;
        RECT 42.200 91.800 42.600 92.200 ;
        RECT 42.200 88.200 42.500 91.800 ;
        RECT 43.000 90.200 43.300 94.800 ;
        RECT 43.000 89.800 43.400 90.200 ;
        RECT 43.800 89.200 44.100 95.800 ;
        RECT 45.400 95.200 45.700 95.800 ;
        RECT 47.800 95.200 48.100 97.800 ;
        RECT 49.400 96.800 49.800 97.200 ;
        RECT 49.400 95.200 49.700 96.800 ;
        RECT 45.400 94.800 45.800 95.200 ;
        RECT 47.800 94.800 48.200 95.200 ;
        RECT 49.400 94.800 49.800 95.200 ;
        RECT 44.600 93.800 45.000 94.200 ;
        RECT 45.400 94.100 45.800 94.200 ;
        RECT 46.200 94.100 46.600 94.200 ;
        RECT 45.400 93.800 46.600 94.100 ;
        RECT 47.000 94.100 47.400 94.200 ;
        RECT 48.600 94.100 49.000 94.200 ;
        RECT 47.000 93.800 49.000 94.100 ;
        RECT 51.000 93.800 51.400 94.200 ;
        RECT 44.600 92.200 44.900 93.800 ;
        RECT 44.600 91.800 45.000 92.200 ;
        RECT 43.800 88.800 44.200 89.200 ;
        RECT 45.400 88.800 45.800 89.200 ;
        RECT 49.400 89.100 49.800 89.200 ;
        RECT 50.200 89.100 50.600 89.200 ;
        RECT 49.400 88.800 50.600 89.100 ;
        RECT 42.200 87.800 42.600 88.200 ;
        RECT 43.800 87.800 44.200 88.200 ;
        RECT 41.400 81.800 41.800 82.200 ;
        RECT 42.200 80.200 42.500 87.800 ;
        RECT 43.800 87.200 44.100 87.800 ;
        RECT 45.400 87.200 45.700 88.800 ;
        RECT 43.800 86.800 44.200 87.200 ;
        RECT 45.400 86.800 45.800 87.200 ;
        RECT 45.400 86.200 45.700 86.800 ;
        RECT 45.400 85.800 45.800 86.200 ;
        RECT 42.200 79.800 42.600 80.200 ;
        RECT 45.400 79.200 45.700 85.800 ;
        RECT 51.000 82.100 51.300 93.800 ;
        RECT 51.800 83.100 52.200 88.900 ;
        RECT 52.600 82.200 52.900 105.800 ;
        RECT 56.600 104.200 56.900 105.800 ;
        RECT 56.600 103.800 57.000 104.200 ;
        RECT 55.800 102.800 56.200 103.200 ;
        RECT 55.800 96.200 56.100 102.800 ;
        RECT 58.200 102.200 58.500 105.800 ;
        RECT 58.200 101.800 58.600 102.200 ;
        RECT 58.200 97.200 58.500 101.800 ;
        RECT 60.600 101.200 60.900 106.800 ;
        RECT 60.600 100.800 61.000 101.200 ;
        RECT 58.200 96.800 58.600 97.200 ;
        RECT 55.800 95.800 56.200 96.200 ;
        RECT 57.400 96.100 57.800 96.200 ;
        RECT 57.400 95.800 58.500 96.100 ;
        RECT 58.200 95.200 58.500 95.800 ;
        RECT 55.000 95.100 55.400 95.200 ;
        RECT 55.800 95.100 56.200 95.200 ;
        RECT 55.000 94.800 56.200 95.100 ;
        RECT 57.400 94.800 57.800 95.200 ;
        RECT 58.200 94.800 58.600 95.200 ;
        RECT 57.400 94.200 57.700 94.800 ;
        RECT 53.400 93.800 53.800 94.200 ;
        RECT 57.400 93.800 57.800 94.200 ;
        RECT 58.200 94.100 58.600 94.200 ;
        RECT 59.000 94.100 59.400 94.200 ;
        RECT 58.200 93.800 59.400 94.100 ;
        RECT 59.800 93.800 60.200 94.200 ;
        RECT 53.400 93.200 53.700 93.800 ;
        RECT 53.400 92.800 53.800 93.200 ;
        RECT 59.800 92.200 60.100 93.800 ;
        RECT 61.400 93.200 61.700 106.800 ;
        RECT 63.800 106.200 64.100 112.800 ;
        RECT 64.600 110.200 64.900 115.800 ;
        RECT 65.400 112.200 65.700 123.800 ;
        RECT 67.800 123.200 68.100 124.800 ;
        RECT 67.800 122.800 68.200 123.200 ;
        RECT 65.400 111.800 65.800 112.200 ;
        RECT 67.000 112.100 67.400 117.900 ;
        RECT 67.800 115.200 68.100 122.800 ;
        RECT 68.600 121.200 68.900 124.800 ;
        RECT 74.200 124.200 74.500 133.800 ;
        RECT 75.800 132.800 76.200 133.200 ;
        RECT 75.800 132.200 76.100 132.800 ;
        RECT 75.000 131.800 75.400 132.200 ;
        RECT 75.800 131.800 76.200 132.200 ;
        RECT 75.000 130.100 75.300 131.800 ;
        RECT 76.600 131.200 76.900 133.800 ;
        RECT 81.400 132.200 81.700 133.800 ;
        RECT 80.600 131.800 81.000 132.200 ;
        RECT 81.400 131.800 81.800 132.200 ;
        RECT 82.200 131.800 82.600 132.200 ;
        RECT 84.600 132.100 85.000 137.900 ;
        RECT 76.600 130.800 77.000 131.200 ;
        RECT 78.200 130.800 78.600 131.200 ;
        RECT 75.000 129.800 76.100 130.100 ;
        RECT 74.200 123.800 74.600 124.200 ;
        RECT 75.000 123.100 75.400 128.900 ;
        RECT 75.800 125.200 76.100 129.800 ;
        RECT 78.200 127.200 78.500 130.800 ;
        RECT 78.200 126.800 78.600 127.200 ;
        RECT 76.600 126.100 77.000 126.200 ;
        RECT 77.400 126.100 77.800 126.200 ;
        RECT 76.600 125.800 77.800 126.100 ;
        RECT 75.800 124.800 76.200 125.200 ;
        RECT 78.200 123.200 78.500 126.800 ;
        RECT 78.200 122.800 78.600 123.200 ;
        RECT 79.000 122.800 79.400 123.200 ;
        RECT 79.800 123.100 80.200 128.900 ;
        RECT 80.600 126.200 80.900 131.800 ;
        RECT 82.200 130.200 82.500 131.800 ;
        RECT 82.200 129.800 82.600 130.200 ;
        RECT 85.400 128.200 85.700 141.800 ;
        RECT 80.600 125.800 81.000 126.200 ;
        RECT 81.400 125.100 81.800 127.900 ;
        RECT 83.800 127.800 84.200 128.200 ;
        RECT 85.400 127.800 85.800 128.200 ;
        RECT 83.800 126.200 84.100 127.800 ;
        RECT 86.200 127.200 86.500 146.800 ;
        RECT 87.000 145.800 87.400 146.200 ;
        RECT 87.000 143.200 87.300 145.800 ;
        RECT 89.400 144.800 89.800 145.200 ;
        RECT 89.400 143.200 89.700 144.800 ;
        RECT 87.000 142.800 87.400 143.200 ;
        RECT 89.400 142.800 89.800 143.200 ;
        RECT 94.200 143.100 94.600 148.900 ;
        RECT 95.000 148.800 95.400 149.200 ;
        RECT 95.000 146.200 95.300 148.800 ;
        RECT 95.800 146.800 96.200 147.200 ;
        RECT 95.800 146.200 96.100 146.800 ;
        RECT 95.000 145.800 95.400 146.200 ;
        RECT 95.800 145.800 96.200 146.200 ;
        RECT 99.000 143.100 99.400 148.900 ;
        RECT 99.800 146.200 100.100 151.800 ;
        RECT 99.800 145.800 100.200 146.200 ;
        RECT 100.600 145.100 101.000 147.900 ;
        RECT 101.400 146.800 101.800 147.200 ;
        RECT 104.600 146.800 105.000 147.200 ;
        RECT 91.800 141.800 92.200 142.200 ;
        RECT 88.600 135.800 89.000 136.200 ;
        RECT 88.600 135.100 88.900 135.800 ;
        RECT 88.600 134.700 89.000 135.100 ;
        RECT 87.000 133.800 87.400 134.200 ;
        RECT 87.000 131.200 87.300 133.800 ;
        RECT 89.400 132.100 89.800 137.900 ;
        RECT 91.800 137.200 92.100 141.800 ;
        RECT 101.400 137.200 101.700 146.800 ;
        RECT 104.600 146.200 104.900 146.800 ;
        RECT 105.400 146.200 105.700 166.800 ;
        RECT 107.000 166.200 107.300 166.800 ;
        RECT 114.200 166.200 114.500 166.800 ;
        RECT 115.800 166.200 116.100 166.800 ;
        RECT 119.000 166.200 119.300 171.800 ;
        RECT 121.400 168.200 121.700 172.800 ;
        RECT 122.200 172.100 122.600 172.200 ;
        RECT 123.000 172.100 123.400 172.200 ;
        RECT 122.200 171.800 123.400 172.100 ;
        RECT 125.400 168.200 125.700 172.800 ;
        RECT 127.000 171.800 127.400 172.200 ;
        RECT 128.600 171.800 129.000 172.200 ;
        RECT 135.800 172.100 136.200 178.900 ;
        RECT 136.600 172.100 137.000 178.900 ;
        RECT 137.400 172.100 137.800 178.900 ;
        RECT 138.200 172.100 138.600 177.900 ;
        RECT 139.000 173.800 139.400 174.200 ;
        RECT 139.000 173.200 139.300 173.800 ;
        RECT 139.000 172.800 139.400 173.200 ;
        RECT 139.800 172.100 140.200 177.900 ;
        RECT 140.600 173.800 141.000 174.200 ;
        RECT 126.200 169.800 126.600 170.200 ;
        RECT 126.200 169.200 126.500 169.800 ;
        RECT 126.200 168.800 126.600 169.200 ;
        RECT 121.400 167.800 121.800 168.200 ;
        RECT 123.800 168.100 124.200 168.200 ;
        RECT 124.600 168.100 125.000 168.200 ;
        RECT 123.800 167.800 125.000 168.100 ;
        RECT 125.400 167.800 125.800 168.200 ;
        RECT 123.800 166.200 124.100 167.800 ;
        RECT 124.600 166.800 125.000 167.200 ;
        RECT 125.400 166.800 125.800 167.200 ;
        RECT 107.000 165.800 107.400 166.200 ;
        RECT 109.400 165.800 109.800 166.200 ;
        RECT 111.000 166.100 111.400 166.200 ;
        RECT 111.800 166.100 112.200 166.200 ;
        RECT 111.000 165.800 112.200 166.100 ;
        RECT 114.200 165.800 114.600 166.200 ;
        RECT 115.800 165.800 116.200 166.200 ;
        RECT 118.200 166.100 118.600 166.200 ;
        RECT 119.000 166.100 119.400 166.200 ;
        RECT 118.200 165.800 119.400 166.100 ;
        RECT 120.600 165.800 121.000 166.200 ;
        RECT 121.400 165.800 121.800 166.200 ;
        RECT 123.800 165.800 124.200 166.200 ;
        RECT 106.200 164.800 106.600 165.200 ;
        RECT 107.000 164.800 107.400 165.200 ;
        RECT 108.600 164.800 109.000 165.200 ;
        RECT 106.200 164.200 106.500 164.800 ;
        RECT 106.200 163.800 106.600 164.200 ;
        RECT 107.000 163.200 107.300 164.800 ;
        RECT 108.600 164.200 108.900 164.800 ;
        RECT 108.600 163.800 109.000 164.200 ;
        RECT 107.000 162.800 107.400 163.200 ;
        RECT 108.600 156.800 109.000 157.200 ;
        RECT 108.600 156.200 108.900 156.800 ;
        RECT 108.600 155.800 109.000 156.200 ;
        RECT 106.200 155.100 106.600 155.200 ;
        RECT 107.000 155.100 107.400 155.200 ;
        RECT 106.200 154.800 107.400 155.100 ;
        RECT 107.000 153.800 107.400 154.200 ;
        RECT 107.000 151.200 107.300 153.800 ;
        RECT 109.400 152.200 109.700 165.800 ;
        RECT 111.800 165.100 112.200 165.200 ;
        RECT 112.600 165.100 113.000 165.200 ;
        RECT 111.800 164.800 113.000 165.100 ;
        RECT 112.600 158.200 112.900 164.800 ;
        RECT 112.600 157.800 113.000 158.200 ;
        RECT 114.200 157.200 114.500 165.800 ;
        RECT 120.600 165.200 120.900 165.800 ;
        RECT 121.400 165.200 121.700 165.800 ;
        RECT 124.600 165.200 124.900 166.800 ;
        RECT 125.400 166.200 125.700 166.800 ;
        RECT 125.400 165.800 125.800 166.200 ;
        RECT 115.000 164.800 115.400 165.200 ;
        RECT 120.600 164.800 121.000 165.200 ;
        RECT 121.400 164.800 121.800 165.200 ;
        RECT 124.600 164.800 125.000 165.200 ;
        RECT 125.400 165.100 125.800 165.200 ;
        RECT 126.200 165.100 126.600 165.200 ;
        RECT 125.400 164.800 126.600 165.100 ;
        RECT 115.000 162.200 115.300 164.800 ;
        RECT 120.600 164.200 120.900 164.800 ;
        RECT 116.600 164.100 117.000 164.200 ;
        RECT 117.400 164.100 117.800 164.200 ;
        RECT 116.600 163.800 117.800 164.100 ;
        RECT 120.600 163.800 121.000 164.200 ;
        RECT 116.600 163.200 116.900 163.800 ;
        RECT 116.600 162.800 117.000 163.200 ;
        RECT 115.000 161.800 115.400 162.200 ;
        RECT 115.800 161.800 116.200 162.200 ;
        RECT 115.000 157.200 115.300 161.800 ;
        RECT 114.200 156.800 114.600 157.200 ;
        RECT 115.000 156.800 115.400 157.200 ;
        RECT 111.000 154.800 111.400 155.200 ;
        RECT 111.800 155.100 112.200 155.200 ;
        RECT 112.600 155.100 113.000 155.200 ;
        RECT 111.800 154.800 113.000 155.100 ;
        RECT 110.200 153.800 110.600 154.200 ;
        RECT 110.200 153.200 110.500 153.800 ;
        RECT 110.200 152.800 110.600 153.200 ;
        RECT 111.000 152.200 111.300 154.800 ;
        RECT 113.400 153.800 113.800 154.200 ;
        RECT 113.400 153.200 113.700 153.800 ;
        RECT 113.400 152.800 113.800 153.200 ;
        RECT 109.400 151.800 109.800 152.200 ;
        RECT 111.000 151.800 111.400 152.200 ;
        RECT 107.000 150.800 107.400 151.200 ;
        RECT 107.000 146.200 107.300 150.800 ;
        RECT 109.400 146.200 109.700 151.800 ;
        RECT 111.800 149.800 112.200 150.200 ;
        RECT 111.800 147.200 112.100 149.800 ;
        RECT 111.800 146.800 112.200 147.200 ;
        RECT 113.400 147.100 113.800 147.200 ;
        RECT 114.200 147.100 114.500 156.800 ;
        RECT 115.800 156.200 116.100 161.800 ;
        RECT 116.600 157.800 117.000 158.200 ;
        RECT 116.600 156.200 116.900 157.800 ;
        RECT 117.400 156.800 117.800 157.200 ;
        RECT 115.800 155.800 116.200 156.200 ;
        RECT 116.600 155.800 117.000 156.200 ;
        RECT 115.000 154.800 115.400 155.200 ;
        RECT 115.000 154.200 115.300 154.800 ;
        RECT 115.000 153.800 115.400 154.200 ;
        RECT 113.400 146.800 114.500 147.100 ;
        RECT 103.800 146.100 104.200 146.200 ;
        RECT 104.600 146.100 105.000 146.200 ;
        RECT 103.800 145.800 105.000 146.100 ;
        RECT 105.400 145.800 105.800 146.200 ;
        RECT 106.200 145.800 106.600 146.200 ;
        RECT 107.000 145.800 107.400 146.200 ;
        RECT 109.400 145.800 109.800 146.200 ;
        RECT 106.200 145.200 106.500 145.800 ;
        RECT 111.800 145.200 112.100 146.800 ;
        RECT 114.200 146.100 114.500 146.800 ;
        RECT 115.000 146.100 115.400 146.200 ;
        RECT 114.200 145.800 115.400 146.100 ;
        RECT 117.400 145.200 117.700 156.800 ;
        RECT 119.000 155.800 119.400 156.200 ;
        RECT 119.000 155.200 119.300 155.800 ;
        RECT 119.000 154.800 119.400 155.200 ;
        RECT 119.000 152.200 119.300 154.800 ;
        RECT 119.800 153.800 120.200 154.200 ;
        RECT 118.200 151.800 118.600 152.200 ;
        RECT 119.000 151.800 119.400 152.200 ;
        RECT 118.200 147.200 118.500 151.800 ;
        RECT 119.800 151.200 120.100 153.800 ;
        RECT 119.800 150.800 120.200 151.200 ;
        RECT 120.600 148.200 120.900 163.800 ;
        RECT 123.000 161.800 123.400 162.200 ;
        RECT 123.000 161.200 123.300 161.800 ;
        RECT 123.000 160.800 123.400 161.200 ;
        RECT 124.600 159.200 124.900 164.800 ;
        RECT 121.400 158.800 121.800 159.200 ;
        RECT 124.600 158.800 125.000 159.200 ;
        RECT 121.400 156.200 121.700 158.800 ;
        RECT 121.400 155.800 121.800 156.200 ;
        RECT 124.600 155.800 125.000 156.200 ;
        RECT 121.400 154.200 121.700 155.800 ;
        RECT 121.400 154.100 121.800 154.200 ;
        RECT 122.200 154.100 122.600 154.200 ;
        RECT 121.400 153.800 122.600 154.100 ;
        RECT 121.400 151.800 121.800 152.200 ;
        RECT 123.000 152.100 123.400 152.200 ;
        RECT 123.800 152.100 124.200 152.200 ;
        RECT 123.000 151.800 124.200 152.100 ;
        RECT 121.400 148.200 121.700 151.800 ;
        RECT 123.800 150.800 124.200 151.200 ;
        RECT 119.000 147.800 119.400 148.200 ;
        RECT 120.600 147.800 121.000 148.200 ;
        RECT 121.400 147.800 121.800 148.200 ;
        RECT 118.200 146.800 118.600 147.200 ;
        RECT 118.200 145.800 118.600 146.200 ;
        RECT 102.200 145.100 102.600 145.200 ;
        RECT 103.000 145.100 103.400 145.200 ;
        RECT 102.200 144.800 103.400 145.100 ;
        RECT 106.200 144.800 106.600 145.200 ;
        RECT 111.800 144.800 112.200 145.200 ;
        RECT 114.200 145.100 114.600 145.200 ;
        RECT 115.000 145.100 115.400 145.200 ;
        RECT 114.200 144.800 115.400 145.100 ;
        RECT 117.400 144.800 117.800 145.200 ;
        RECT 117.400 144.200 117.700 144.800 ;
        RECT 103.800 143.800 104.200 144.200 ;
        RECT 107.000 143.800 107.400 144.200 ;
        RECT 107.800 143.800 108.200 144.200 ;
        RECT 110.200 143.800 110.600 144.200 ;
        RECT 115.800 143.800 116.200 144.200 ;
        RECT 117.400 143.800 117.800 144.200 ;
        RECT 103.800 140.200 104.100 143.800 ;
        RECT 107.000 143.200 107.300 143.800 ;
        RECT 107.000 142.800 107.400 143.200 ;
        RECT 107.800 140.200 108.100 143.800 ;
        RECT 109.400 141.800 109.800 142.200 ;
        RECT 103.800 139.800 104.200 140.200 ;
        RECT 107.800 139.800 108.200 140.200 ;
        RECT 109.400 139.200 109.700 141.800 ;
        RECT 109.400 138.800 109.800 139.200 ;
        RECT 103.800 137.800 104.200 138.200 ;
        RECT 105.400 137.800 105.800 138.200 ;
        RECT 91.800 136.800 92.200 137.200 ;
        RECT 101.400 136.800 101.800 137.200 ;
        RECT 91.000 133.100 91.400 135.900 ;
        RECT 93.400 135.800 93.800 136.200 ;
        RECT 102.200 135.800 102.600 136.200 ;
        RECT 93.400 134.200 93.700 135.800 ;
        RECT 102.200 135.200 102.500 135.800 ;
        RECT 94.200 134.800 94.600 135.200 ;
        RECT 95.800 134.800 96.200 135.200 ;
        RECT 102.200 134.800 102.600 135.200 ;
        RECT 94.200 134.200 94.500 134.800 ;
        RECT 91.800 133.800 92.200 134.200 ;
        RECT 93.400 133.800 93.800 134.200 ;
        RECT 94.200 133.800 94.600 134.200 ;
        RECT 87.000 130.800 87.400 131.200 ;
        RECT 91.800 130.200 92.100 133.800 ;
        RECT 92.600 130.800 93.000 131.200 ;
        RECT 87.000 129.800 87.400 130.200 ;
        RECT 91.800 129.800 92.200 130.200 ;
        RECT 87.000 128.200 87.300 129.800 ;
        RECT 89.400 129.100 89.800 129.200 ;
        RECT 90.200 129.100 90.600 129.200 ;
        RECT 89.400 128.800 90.600 129.100 ;
        RECT 87.000 127.800 87.400 128.200 ;
        RECT 87.800 128.100 88.200 128.200 ;
        RECT 88.600 128.100 89.000 128.200 ;
        RECT 87.800 127.800 89.000 128.100 ;
        RECT 84.600 126.800 85.000 127.200 ;
        RECT 86.200 126.800 86.600 127.200 ;
        RECT 83.800 125.800 84.200 126.200 ;
        RECT 82.200 125.100 82.600 125.200 ;
        RECT 83.000 125.100 83.400 125.200 ;
        RECT 82.200 124.800 83.400 125.100 ;
        RECT 84.600 124.200 84.900 126.800 ;
        RECT 85.400 126.100 85.800 126.200 ;
        RECT 86.200 126.100 86.600 126.200 ;
        RECT 85.400 125.800 86.600 126.100 ;
        RECT 86.200 124.200 86.500 125.800 ;
        RECT 84.600 123.800 85.000 124.200 ;
        RECT 86.200 123.800 86.600 124.200 ;
        RECT 91.800 123.100 92.200 128.900 ;
        RECT 92.600 126.200 92.900 130.800 ;
        RECT 92.600 126.100 93.000 126.200 ;
        RECT 94.200 126.100 94.600 126.200 ;
        RECT 95.000 126.100 95.400 126.200 ;
        RECT 92.600 125.800 93.700 126.100 ;
        RECT 94.200 125.800 95.400 126.100 ;
        RECT 72.600 121.800 73.000 122.200 ;
        RECT 75.000 121.800 75.400 122.200 ;
        RECT 68.600 120.800 69.000 121.200 ;
        RECT 67.800 114.800 68.200 115.200 ;
        RECT 70.200 114.800 70.600 115.200 ;
        RECT 67.800 111.800 68.200 112.200 ;
        RECT 64.600 109.800 65.000 110.200 ;
        RECT 67.000 109.800 67.400 110.200 ;
        RECT 67.000 109.200 67.300 109.800 ;
        RECT 64.600 108.800 65.000 109.200 ;
        RECT 67.000 108.800 67.400 109.200 ;
        RECT 64.600 108.200 64.900 108.800 ;
        RECT 64.600 107.800 65.000 108.200 ;
        RECT 66.200 108.100 66.600 108.200 ;
        RECT 66.200 107.800 67.300 108.100 ;
        RECT 67.000 107.200 67.300 107.800 ;
        RECT 67.800 107.200 68.100 111.800 ;
        RECT 70.200 111.200 70.500 114.800 ;
        RECT 71.800 112.100 72.200 117.900 ;
        RECT 70.200 110.800 70.600 111.200 ;
        RECT 71.800 109.800 72.200 110.200 ;
        RECT 71.800 109.200 72.100 109.800 ;
        RECT 70.200 108.800 70.600 109.200 ;
        RECT 71.800 108.800 72.200 109.200 ;
        RECT 69.400 107.800 69.800 108.200 ;
        RECT 69.400 107.200 69.700 107.800 ;
        RECT 67.000 106.800 67.400 107.200 ;
        RECT 67.800 106.800 68.200 107.200 ;
        RECT 69.400 106.800 69.800 107.200 ;
        RECT 63.800 105.800 64.200 106.200 ;
        RECT 65.400 101.800 65.800 102.200 ;
        RECT 62.200 99.800 62.600 100.200 ;
        RECT 64.600 99.800 65.000 100.200 ;
        RECT 62.200 99.200 62.500 99.800 ;
        RECT 62.200 98.800 62.600 99.200 ;
        RECT 64.600 95.200 64.900 99.800 ;
        RECT 65.400 97.200 65.700 101.800 ;
        RECT 67.000 99.200 67.300 106.800 ;
        RECT 70.200 106.200 70.500 108.800 ;
        RECT 71.800 107.800 72.200 108.200 ;
        RECT 72.600 108.100 72.900 121.800 ;
        RECT 75.000 119.200 75.300 121.800 ;
        RECT 75.000 118.800 75.400 119.200 ;
        RECT 73.400 113.100 73.800 115.900 ;
        RECT 76.600 115.100 77.000 115.200 ;
        RECT 77.400 115.100 77.800 115.200 ;
        RECT 76.600 114.800 77.800 115.100 ;
        RECT 74.200 113.800 74.600 114.200 ;
        RECT 73.400 108.100 73.800 108.200 ;
        RECT 72.600 107.800 73.800 108.100 ;
        RECT 71.800 106.200 72.100 107.800 ;
        RECT 72.600 106.800 73.000 107.200 ;
        RECT 72.600 106.200 72.900 106.800 ;
        RECT 68.600 106.100 69.000 106.200 ;
        RECT 69.400 106.100 69.800 106.200 ;
        RECT 68.600 105.800 69.800 106.100 ;
        RECT 70.200 105.800 70.600 106.200 ;
        RECT 71.800 105.800 72.200 106.200 ;
        RECT 72.600 105.800 73.000 106.200 ;
        RECT 67.800 104.800 68.200 105.200 ;
        RECT 67.000 98.800 67.400 99.200 ;
        RECT 65.400 96.800 65.800 97.200 ;
        RECT 64.600 94.800 65.000 95.200 ;
        RECT 65.400 95.100 65.800 95.200 ;
        RECT 66.200 95.100 66.600 95.200 ;
        RECT 65.400 94.800 66.600 95.100 ;
        RECT 63.800 94.100 64.200 94.200 ;
        RECT 64.600 94.100 65.000 94.200 ;
        RECT 63.800 93.800 65.000 94.100 ;
        RECT 61.400 92.800 61.800 93.200 ;
        RECT 59.800 91.800 60.200 92.200 ;
        RECT 61.400 91.200 61.700 92.800 ;
        RECT 64.600 91.800 65.000 92.200 ;
        RECT 55.800 90.800 56.200 91.200 ;
        RECT 61.400 90.800 61.800 91.200 ;
        RECT 55.800 88.200 56.100 90.800 ;
        RECT 55.800 87.800 56.200 88.200 ;
        RECT 55.000 86.200 55.400 86.300 ;
        RECT 55.800 86.200 56.200 86.300 ;
        RECT 55.000 85.900 56.200 86.200 ;
        RECT 56.600 83.100 57.000 88.900 ;
        RECT 59.000 88.800 59.400 89.200 ;
        RECT 63.800 88.800 64.200 89.200 ;
        RECT 58.200 85.100 58.600 87.900 ;
        RECT 59.000 87.200 59.300 88.800 ;
        RECT 63.000 87.800 63.400 88.200 ;
        RECT 59.000 86.800 59.400 87.200 ;
        RECT 60.600 86.800 61.000 87.200 ;
        RECT 60.600 86.200 60.900 86.800 ;
        RECT 63.000 86.200 63.300 87.800 ;
        RECT 63.800 87.200 64.100 88.800 ;
        RECT 63.800 86.800 64.200 87.200 ;
        RECT 64.600 86.200 64.900 91.800 ;
        RECT 67.000 90.800 67.400 91.200 ;
        RECT 66.200 89.800 66.600 90.200 ;
        RECT 66.200 89.200 66.500 89.800 ;
        RECT 66.200 88.800 66.600 89.200 ;
        RECT 67.000 86.200 67.300 90.800 ;
        RECT 67.800 89.200 68.100 104.800 ;
        RECT 69.400 103.800 69.800 104.200 ;
        RECT 69.400 99.200 69.700 103.800 ;
        RECT 71.800 100.200 72.100 105.800 ;
        RECT 74.200 103.100 74.500 113.800 ;
        RECT 76.600 113.200 76.900 114.800 ;
        RECT 76.600 112.800 77.000 113.200 ;
        RECT 75.000 106.800 75.400 107.200 ;
        RECT 75.000 106.200 75.300 106.800 ;
        RECT 75.000 105.800 75.400 106.200 ;
        RECT 75.800 105.100 76.200 107.900 ;
        RECT 77.400 103.100 77.800 108.900 ;
        RECT 78.200 108.200 78.500 122.800 ;
        RECT 79.000 119.200 79.300 122.800 ;
        RECT 83.800 121.800 84.200 122.200 ;
        RECT 86.200 121.800 86.600 122.200 ;
        RECT 83.800 120.100 84.100 121.800 ;
        RECT 83.800 119.800 84.900 120.100 ;
        RECT 79.000 118.800 79.400 119.200 ;
        RECT 83.800 118.800 84.200 119.200 ;
        RECT 79.800 114.800 80.200 115.200 ;
        RECT 79.800 114.200 80.100 114.800 ;
        RECT 79.800 113.800 80.200 114.200 ;
        RECT 83.000 113.800 83.400 114.200 ;
        RECT 79.000 111.800 79.400 112.200 ;
        RECT 82.200 111.800 82.600 112.200 ;
        RECT 78.200 107.800 78.600 108.200 ;
        RECT 73.400 102.800 74.500 103.100 ;
        RECT 73.400 102.200 73.700 102.800 ;
        RECT 73.400 101.800 73.800 102.200 ;
        RECT 74.200 101.800 74.600 102.200 ;
        RECT 71.800 99.800 72.200 100.200 ;
        RECT 69.400 98.800 69.800 99.200 ;
        RECT 71.800 98.800 72.200 99.200 ;
        RECT 71.800 94.200 72.100 98.800 ;
        RECT 73.400 95.200 73.700 101.800 ;
        RECT 74.200 98.200 74.500 101.800 ;
        RECT 75.800 100.800 76.200 101.200 ;
        RECT 74.200 97.800 74.600 98.200 ;
        RECT 75.800 95.200 76.100 100.800 ;
        RECT 78.200 98.800 78.600 99.200 ;
        RECT 76.600 96.800 77.000 97.200 ;
        RECT 76.600 96.200 76.900 96.800 ;
        RECT 76.600 95.800 77.000 96.200 ;
        RECT 78.200 95.200 78.500 98.800 ;
        RECT 79.000 97.200 79.300 111.800 ;
        RECT 82.200 110.200 82.500 111.800 ;
        RECT 82.200 109.800 82.600 110.200 ;
        RECT 83.000 109.200 83.300 113.800 ;
        RECT 83.800 113.200 84.100 118.800 ;
        RECT 84.600 114.100 84.900 119.800 ;
        RECT 85.400 118.100 85.800 118.200 ;
        RECT 86.200 118.100 86.500 121.800 ;
        RECT 85.400 117.800 86.500 118.100 ;
        RECT 87.000 117.800 87.400 118.200 ;
        RECT 86.200 115.800 86.600 116.200 ;
        RECT 86.200 115.200 86.500 115.800 ;
        RECT 87.000 115.200 87.300 117.800 ;
        RECT 91.800 116.800 92.200 117.200 ;
        RECT 91.800 116.200 92.100 116.800 ;
        RECT 87.800 115.800 88.200 116.200 ;
        RECT 91.800 115.800 92.200 116.200 ;
        RECT 87.800 115.200 88.100 115.800 ;
        RECT 86.200 114.800 86.600 115.200 ;
        RECT 87.000 114.800 87.400 115.200 ;
        RECT 87.800 114.800 88.200 115.200 ;
        RECT 86.200 114.200 86.500 114.800 ;
        RECT 85.400 114.100 85.800 114.200 ;
        RECT 84.600 113.800 85.800 114.100 ;
        RECT 86.200 113.800 86.600 114.200 ;
        RECT 88.600 113.800 89.000 114.200 ;
        RECT 89.400 113.800 89.800 114.200 ;
        RECT 90.200 113.800 90.600 114.200 ;
        RECT 83.800 112.800 84.200 113.200 ;
        RECT 79.800 107.800 80.200 108.200 ;
        RECT 79.800 106.200 80.100 107.800 ;
        RECT 79.800 105.800 80.200 106.200 ;
        RECT 82.200 103.100 82.600 108.900 ;
        RECT 83.000 108.800 83.400 109.200 ;
        RECT 80.600 100.800 81.000 101.200 ;
        RECT 79.000 96.800 79.400 97.200 ;
        RECT 79.000 96.100 79.300 96.800 ;
        RECT 79.800 96.100 80.200 96.200 ;
        RECT 79.000 95.800 80.200 96.100 ;
        RECT 73.400 94.800 73.800 95.200 ;
        RECT 74.200 94.800 74.600 95.200 ;
        RECT 75.000 94.800 75.400 95.200 ;
        RECT 75.800 94.800 76.200 95.200 ;
        RECT 78.200 95.100 78.600 95.200 ;
        RECT 79.000 95.100 79.400 95.200 ;
        RECT 78.200 94.800 79.400 95.100 ;
        RECT 74.200 94.200 74.500 94.800 ;
        RECT 71.800 93.800 72.200 94.200 ;
        RECT 72.600 93.800 73.000 94.200 ;
        RECT 74.200 93.800 74.600 94.200 ;
        RECT 68.600 92.100 69.000 92.200 ;
        RECT 69.400 92.100 69.800 92.200 ;
        RECT 68.600 91.800 69.800 92.100 ;
        RECT 71.800 89.200 72.100 93.800 ;
        RECT 72.600 91.200 72.900 93.800 ;
        RECT 73.400 91.800 73.800 92.200 ;
        RECT 72.600 90.800 73.000 91.200 ;
        RECT 67.800 88.800 68.200 89.200 ;
        RECT 71.800 88.800 72.200 89.200 ;
        RECT 73.400 87.200 73.700 91.800 ;
        RECT 75.000 89.200 75.300 94.800 ;
        RECT 75.800 93.800 76.200 94.200 ;
        RECT 78.200 94.100 78.600 94.200 ;
        RECT 79.000 94.100 79.400 94.200 ;
        RECT 78.200 93.800 79.400 94.100 ;
        RECT 75.800 93.200 76.100 93.800 ;
        RECT 75.800 92.800 76.200 93.200 ;
        RECT 74.200 88.800 74.600 89.200 ;
        RECT 75.000 88.800 75.400 89.200 ;
        RECT 74.200 88.200 74.500 88.800 ;
        RECT 74.200 87.800 74.600 88.200 ;
        RECT 80.600 87.200 80.900 100.800 ;
        RECT 81.400 98.800 81.800 99.200 ;
        RECT 81.400 98.200 81.700 98.800 ;
        RECT 81.400 97.800 81.800 98.200 ;
        RECT 83.000 96.800 83.400 97.200 ;
        RECT 83.000 96.200 83.300 96.800 ;
        RECT 83.000 95.800 83.400 96.200 ;
        RECT 83.000 95.100 83.400 95.200 ;
        RECT 83.800 95.100 84.100 112.800 ;
        RECT 84.600 109.100 85.000 109.200 ;
        RECT 85.400 109.100 85.800 109.200 ;
        RECT 84.600 108.800 85.800 109.100 ;
        RECT 87.800 108.800 88.200 109.200 ;
        RECT 85.400 106.800 85.800 107.200 ;
        RECT 87.000 106.800 87.400 107.200 ;
        RECT 85.400 106.200 85.700 106.800 ;
        RECT 87.000 106.200 87.300 106.800 ;
        RECT 87.800 106.200 88.100 108.800 ;
        RECT 88.600 108.200 88.900 113.800 ;
        RECT 89.400 108.200 89.700 113.800 ;
        RECT 90.200 109.200 90.500 113.800 ;
        RECT 92.600 113.100 93.000 115.900 ;
        RECT 93.400 114.200 93.700 125.800 ;
        RECT 93.400 113.800 93.800 114.200 ;
        RECT 94.200 112.100 94.600 117.900 ;
        RECT 95.800 115.200 96.100 134.800 ;
        RECT 96.600 134.100 97.000 134.200 ;
        RECT 97.400 134.100 97.800 134.200 ;
        RECT 96.600 133.800 97.800 134.100 ;
        RECT 98.200 132.800 98.600 133.200 ;
        RECT 98.200 132.200 98.500 132.800 ;
        RECT 98.200 131.800 98.600 132.200 ;
        RECT 96.600 123.100 97.000 128.900 ;
        RECT 99.000 128.800 99.400 129.200 ;
        RECT 98.200 125.100 98.600 127.900 ;
        RECT 99.000 127.200 99.300 128.800 ;
        RECT 99.000 126.800 99.400 127.200 ;
        RECT 100.600 127.100 101.000 127.200 ;
        RECT 99.800 126.800 101.000 127.100 ;
        RECT 99.800 126.200 100.100 126.800 ;
        RECT 99.800 125.800 100.200 126.200 ;
        RECT 100.600 125.800 101.000 126.200 ;
        RECT 100.600 125.200 100.900 125.800 ;
        RECT 100.600 124.800 101.000 125.200 ;
        RECT 96.600 115.800 97.000 116.200 ;
        RECT 96.600 115.200 96.900 115.800 ;
        RECT 95.800 114.800 96.200 115.200 ;
        RECT 96.600 114.800 97.000 115.200 ;
        RECT 97.400 112.800 97.800 113.200 ;
        RECT 90.200 108.800 90.600 109.200 ;
        RECT 94.200 108.800 94.600 109.200 ;
        RECT 94.200 108.200 94.500 108.800 ;
        RECT 97.400 108.200 97.700 112.800 ;
        RECT 99.000 112.100 99.400 117.900 ;
        RECT 88.600 107.800 89.000 108.200 ;
        RECT 89.400 108.100 89.800 108.200 ;
        RECT 90.200 108.100 90.600 108.200 ;
        RECT 89.400 107.800 90.600 108.100 ;
        RECT 94.200 107.800 94.600 108.200 ;
        RECT 97.400 107.800 97.800 108.200 ;
        RECT 89.400 106.800 89.800 107.200 ;
        RECT 92.600 107.100 93.000 107.200 ;
        RECT 93.400 107.100 93.800 107.200 ;
        RECT 92.600 106.800 93.800 107.100 ;
        RECT 98.200 106.800 98.600 107.200 ;
        RECT 99.800 106.800 100.200 107.200 ;
        RECT 89.400 106.200 89.700 106.800 ;
        RECT 85.400 105.800 85.800 106.200 ;
        RECT 87.000 105.800 87.400 106.200 ;
        RECT 87.800 105.800 88.200 106.200 ;
        RECT 89.400 105.800 89.800 106.200 ;
        RECT 91.800 105.800 92.200 106.200 ;
        RECT 95.800 106.100 96.200 106.200 ;
        RECT 96.600 106.100 97.000 106.200 ;
        RECT 95.800 105.800 97.000 106.100 ;
        RECT 85.400 104.800 85.800 105.200 ;
        RECT 90.200 105.100 90.600 105.200 ;
        RECT 91.000 105.100 91.400 105.200 ;
        RECT 90.200 104.800 91.400 105.100 ;
        RECT 85.400 104.200 85.700 104.800 ;
        RECT 85.400 103.800 85.800 104.200 ;
        RECT 90.200 103.800 90.600 104.200 ;
        RECT 88.600 101.800 89.000 102.200 ;
        RECT 86.200 96.800 86.600 97.200 ;
        RECT 83.000 94.800 84.100 95.100 ;
        RECT 84.600 95.100 85.000 95.200 ;
        RECT 85.400 95.100 85.800 95.200 ;
        RECT 84.600 94.800 85.800 95.100 ;
        RECT 86.200 94.200 86.500 96.800 ;
        RECT 88.600 95.200 88.900 101.800 ;
        RECT 90.200 99.200 90.500 103.800 ;
        RECT 91.000 103.200 91.300 104.800 ;
        RECT 91.800 104.200 92.100 105.800 ;
        RECT 97.400 104.800 97.800 105.200 ;
        RECT 91.800 103.800 92.200 104.200 ;
        RECT 91.000 102.800 91.400 103.200 ;
        RECT 94.200 101.800 94.600 102.200 ;
        RECT 96.600 101.800 97.000 102.200 ;
        RECT 90.200 98.800 90.600 99.200 ;
        RECT 93.400 98.800 93.800 99.200 ;
        RECT 91.800 97.800 92.200 98.200 ;
        RECT 87.000 94.800 87.400 95.200 ;
        RECT 88.600 94.800 89.000 95.200 ;
        RECT 82.200 94.100 82.600 94.200 ;
        RECT 81.400 93.800 82.600 94.100 ;
        RECT 85.400 93.800 85.800 94.200 ;
        RECT 86.200 93.800 86.600 94.200 ;
        RECT 70.200 86.800 70.600 87.200 ;
        RECT 73.400 86.800 73.800 87.200 ;
        RECT 75.000 87.100 75.400 87.200 ;
        RECT 75.800 87.100 76.200 87.200 ;
        RECT 75.000 86.800 76.200 87.100 ;
        RECT 79.800 86.800 80.200 87.200 ;
        RECT 80.600 86.800 81.000 87.200 ;
        RECT 60.600 85.800 61.000 86.200 ;
        RECT 63.000 85.800 63.400 86.200 ;
        RECT 64.600 85.800 65.000 86.200 ;
        RECT 67.000 85.800 67.400 86.200 ;
        RECT 69.400 85.800 69.800 86.200 ;
        RECT 63.000 85.200 63.300 85.800 ;
        RECT 60.600 85.100 61.000 85.200 ;
        RECT 61.400 85.100 61.800 85.200 ;
        RECT 60.600 84.800 61.800 85.100 ;
        RECT 63.000 84.800 63.400 85.200 ;
        RECT 64.600 83.200 64.900 85.800 ;
        RECT 67.800 83.800 68.200 84.200 ;
        RECT 64.600 82.800 65.000 83.200 ;
        RECT 65.400 82.800 65.800 83.200 ;
        RECT 51.000 81.800 52.100 82.100 ;
        RECT 52.600 81.800 53.000 82.200 ;
        RECT 58.200 81.800 58.600 82.200 ;
        RECT 47.800 79.800 48.200 80.200 ;
        RECT 45.400 78.800 45.800 79.200 ;
        RECT 39.000 72.100 39.400 77.900 ;
        RECT 42.200 77.800 42.600 78.200 ;
        RECT 42.200 77.200 42.500 77.800 ;
        RECT 39.800 76.800 40.200 77.200 ;
        RECT 42.200 76.800 42.600 77.200 ;
        RECT 38.200 58.800 38.600 59.200 ;
        RECT 34.200 56.800 34.600 57.200 ;
        RECT 35.000 56.800 35.400 57.200 ;
        RECT 32.600 49.100 33.000 49.200 ;
        RECT 33.400 49.100 33.800 49.200 ;
        RECT 31.000 43.100 31.400 48.900 ;
        RECT 32.600 48.800 33.800 49.100 ;
        RECT 34.200 47.200 34.500 56.800 ;
        RECT 39.800 56.200 40.100 76.800 ;
        RECT 42.200 74.200 42.500 76.800 ;
        RECT 43.800 76.100 44.200 76.200 ;
        RECT 44.600 76.100 45.000 76.200 ;
        RECT 43.800 75.800 45.000 76.100 ;
        RECT 47.800 75.200 48.100 79.800 ;
        RECT 50.200 78.800 50.600 79.200 ;
        RECT 50.200 76.200 50.500 78.800 ;
        RECT 48.600 76.100 49.000 76.200 ;
        RECT 50.200 76.100 50.600 76.200 ;
        RECT 51.000 76.100 51.400 76.200 ;
        RECT 48.600 75.800 49.700 76.100 ;
        RECT 50.200 75.800 51.400 76.100 ;
        RECT 49.400 75.200 49.700 75.800 ;
        RECT 43.800 74.800 44.200 75.200 ;
        RECT 46.200 75.100 46.600 75.200 ;
        RECT 47.000 75.100 47.400 75.200 ;
        RECT 46.200 74.800 47.400 75.100 ;
        RECT 47.800 74.800 48.200 75.200 ;
        RECT 48.600 74.800 49.000 75.200 ;
        RECT 49.400 74.800 49.800 75.200 ;
        RECT 51.000 74.800 51.400 75.200 ;
        RECT 43.800 74.200 44.100 74.800 ;
        RECT 47.800 74.200 48.100 74.800 ;
        RECT 42.200 73.800 42.600 74.200 ;
        RECT 43.800 73.800 44.200 74.200 ;
        RECT 46.200 74.100 46.600 74.200 ;
        RECT 47.000 74.100 47.400 74.200 ;
        RECT 46.200 73.800 47.400 74.100 ;
        RECT 47.800 73.800 48.200 74.200 ;
        RECT 47.800 73.200 48.100 73.800 ;
        RECT 43.800 72.800 44.200 73.200 ;
        RECT 47.800 72.800 48.200 73.200 ;
        RECT 40.600 63.100 41.000 68.900 ;
        RECT 43.800 67.200 44.100 72.800 ;
        RECT 46.200 69.800 46.600 70.200 ;
        RECT 46.200 69.200 46.500 69.800 ;
        RECT 48.600 69.200 48.900 74.800 ;
        RECT 51.000 74.200 51.300 74.800 ;
        RECT 51.000 73.800 51.400 74.200 ;
        RECT 51.800 71.200 52.100 81.800 ;
        RECT 53.400 78.800 53.800 79.200 ;
        RECT 53.400 78.200 53.700 78.800 ;
        RECT 52.600 77.800 53.000 78.200 ;
        RECT 53.400 77.800 53.800 78.200 ;
        RECT 52.600 75.200 52.900 77.800 ;
        RECT 55.000 76.800 55.400 77.200 ;
        RECT 55.000 76.200 55.300 76.800 ;
        RECT 54.200 75.800 54.600 76.200 ;
        RECT 55.000 75.800 55.400 76.200 ;
        RECT 52.600 74.800 53.000 75.200 ;
        RECT 53.400 73.800 53.800 74.200 ;
        RECT 51.800 70.800 52.200 71.200 ;
        RECT 46.200 68.800 46.600 69.200 ;
        RECT 48.600 68.800 49.000 69.200 ;
        RECT 47.800 68.100 48.200 68.200 ;
        RECT 48.600 68.100 49.000 68.200 ;
        RECT 47.800 67.800 49.000 68.100 ;
        RECT 49.400 68.100 49.800 68.200 ;
        RECT 50.200 68.100 50.600 68.200 ;
        RECT 49.400 67.800 50.600 68.100 ;
        RECT 42.200 67.100 42.600 67.200 ;
        RECT 43.000 67.100 43.400 67.200 ;
        RECT 42.200 66.800 43.400 67.100 ;
        RECT 43.800 66.800 44.200 67.200 ;
        RECT 47.000 67.100 47.400 67.200 ;
        RECT 47.800 67.100 48.200 67.200 ;
        RECT 47.000 66.800 48.200 67.100 ;
        RECT 51.000 66.800 51.400 67.200 ;
        RECT 51.800 67.100 52.200 67.200 ;
        RECT 52.600 67.100 53.000 67.200 ;
        RECT 51.800 66.800 53.000 67.100 ;
        RECT 51.000 66.200 51.300 66.800 ;
        RECT 44.600 65.800 45.000 66.200 ;
        RECT 46.200 65.800 46.600 66.200 ;
        RECT 47.000 65.800 47.400 66.200 ;
        RECT 51.000 65.800 51.400 66.200 ;
        RECT 41.400 64.100 41.800 64.200 ;
        RECT 42.200 64.100 42.600 64.200 ;
        RECT 41.400 63.800 42.600 64.100 ;
        RECT 41.400 62.800 41.800 63.200 ;
        RECT 41.400 59.200 41.700 62.800 ;
        RECT 44.600 61.200 44.900 65.800 ;
        RECT 46.200 65.200 46.500 65.800 ;
        RECT 46.200 64.800 46.600 65.200 ;
        RECT 46.200 63.800 46.600 64.200 ;
        RECT 44.600 60.800 45.000 61.200 ;
        RECT 41.400 58.800 41.800 59.200 ;
        RECT 43.000 58.800 43.400 59.200 ;
        RECT 41.400 57.800 41.800 58.200 ;
        RECT 36.600 56.100 37.000 56.200 ;
        RECT 37.400 56.100 37.800 56.200 ;
        RECT 36.600 55.800 37.800 56.100 ;
        RECT 39.800 55.800 40.200 56.200 ;
        RECT 37.400 55.100 37.800 55.200 ;
        RECT 38.200 55.100 38.600 55.200 ;
        RECT 37.400 54.800 38.600 55.100 ;
        RECT 39.000 54.800 39.400 55.200 ;
        RECT 39.000 54.200 39.300 54.800 ;
        RECT 39.800 54.200 40.100 55.800 ;
        RECT 41.400 55.200 41.700 57.800 ;
        RECT 43.000 56.200 43.300 58.800 ;
        RECT 43.000 55.800 43.400 56.200 ;
        RECT 41.400 54.800 41.800 55.200 ;
        RECT 39.000 53.800 39.400 54.200 ;
        RECT 39.800 53.800 40.200 54.200 ;
        RECT 40.600 53.800 41.000 54.200 ;
        RECT 39.000 51.200 39.300 53.800 ;
        RECT 39.000 50.800 39.400 51.200 ;
        RECT 35.000 47.800 35.400 48.200 ;
        RECT 39.000 47.800 39.400 48.200 ;
        RECT 34.200 46.800 34.600 47.200 ;
        RECT 28.600 35.800 29.000 36.200 ;
        RECT 27.000 35.100 27.400 35.200 ;
        RECT 27.800 35.100 28.200 35.200 ;
        RECT 27.000 34.800 28.200 35.100 ;
        RECT 25.400 32.800 25.800 33.200 ;
        RECT 23.000 27.800 23.400 28.200 ;
        RECT 23.000 26.200 23.300 27.800 ;
        RECT 25.400 27.200 25.700 32.800 ;
        RECT 29.400 32.100 29.800 37.900 ;
        RECT 31.800 37.800 32.200 38.200 ;
        RECT 31.800 37.200 32.100 37.800 ;
        RECT 31.800 36.800 32.200 37.200 ;
        RECT 32.600 35.800 33.000 36.200 ;
        RECT 34.200 36.100 34.500 46.800 ;
        RECT 35.000 46.200 35.300 47.800 ;
        RECT 39.000 47.200 39.300 47.800 ;
        RECT 36.600 47.100 37.000 47.200 ;
        RECT 37.400 47.100 37.800 47.200 ;
        RECT 36.600 46.800 37.800 47.100 ;
        RECT 39.000 46.800 39.400 47.200 ;
        RECT 35.000 45.800 35.400 46.200 ;
        RECT 37.400 45.800 37.800 46.200 ;
        RECT 37.400 45.200 37.700 45.800 ;
        RECT 37.400 44.800 37.800 45.200 ;
        RECT 39.800 45.100 40.200 47.900 ;
        RECT 40.600 42.200 40.900 53.800 ;
        RECT 41.400 43.100 41.800 48.900 ;
        RECT 42.200 46.800 42.600 47.200 ;
        RECT 42.200 46.300 42.500 46.800 ;
        RECT 42.200 45.900 42.600 46.300 ;
        RECT 42.200 45.800 42.500 45.900 ;
        RECT 40.600 41.800 41.000 42.200 ;
        RECT 38.200 38.800 38.600 39.200 ;
        RECT 33.400 35.800 34.500 36.100 ;
        RECT 35.800 36.800 36.200 37.200 ;
        RECT 37.400 36.800 37.800 37.200 ;
        RECT 32.600 34.200 32.900 35.800 ;
        RECT 33.400 35.200 33.700 35.800 ;
        RECT 33.400 34.800 33.800 35.200 ;
        RECT 34.200 35.100 34.600 35.200 ;
        RECT 35.000 35.100 35.400 35.200 ;
        RECT 34.200 34.800 35.400 35.100 ;
        RECT 30.200 33.800 30.600 34.200 ;
        RECT 32.600 33.800 33.000 34.200 ;
        RECT 28.600 30.800 29.000 31.200 ;
        RECT 28.600 29.200 28.900 30.800 ;
        RECT 25.400 26.800 25.800 27.200 ;
        RECT 22.200 25.800 22.600 26.200 ;
        RECT 23.000 25.800 23.400 26.200 ;
        RECT 26.200 23.100 26.600 28.900 ;
        RECT 28.600 28.800 29.000 29.200 ;
        RECT 19.000 15.100 19.400 15.200 ;
        RECT 19.800 15.100 20.200 15.200 ;
        RECT 19.000 14.800 20.200 15.100 ;
        RECT 20.600 14.800 21.000 15.200 ;
        RECT 22.200 12.100 22.600 17.900 ;
        RECT 30.200 17.200 30.500 33.800 ;
        RECT 33.400 32.200 33.700 34.800 ;
        RECT 35.800 34.200 36.100 36.800 ;
        RECT 37.400 36.200 37.700 36.800 ;
        RECT 37.400 35.800 37.800 36.200 ;
        RECT 35.800 33.800 36.200 34.200 ;
        RECT 38.200 33.200 38.500 38.800 ;
        RECT 43.000 37.100 43.300 55.800 ;
        RECT 43.800 53.100 44.200 55.900 ;
        RECT 44.600 53.800 45.000 54.200 ;
        RECT 44.600 46.200 44.900 53.800 ;
        RECT 45.400 52.100 45.800 57.900 ;
        RECT 46.200 54.200 46.500 63.800 ;
        RECT 47.000 58.200 47.300 65.800 ;
        RECT 52.600 64.800 53.000 65.200 ;
        RECT 52.600 64.200 52.900 64.800 ;
        RECT 52.600 63.800 53.000 64.200 ;
        RECT 47.000 57.800 47.400 58.200 ;
        RECT 47.000 56.800 47.400 57.200 ;
        RECT 47.000 55.200 47.300 56.800 ;
        RECT 47.000 54.800 47.400 55.200 ;
        RECT 46.200 53.800 46.600 54.200 ;
        RECT 50.200 52.100 50.600 57.900 ;
        RECT 52.600 56.800 53.000 57.200 ;
        RECT 51.000 55.800 51.400 56.200 ;
        RECT 45.400 47.800 45.800 48.200 ;
        RECT 45.400 47.200 45.700 47.800 ;
        RECT 45.400 46.800 45.800 47.200 ;
        RECT 44.600 45.800 45.000 46.200 ;
        RECT 43.800 42.800 44.200 43.200 ;
        RECT 46.200 43.100 46.600 48.900 ;
        RECT 51.000 47.200 51.300 55.800 ;
        RECT 52.600 55.200 52.900 56.800 ;
        RECT 52.600 54.800 53.000 55.200 ;
        RECT 53.400 54.200 53.700 73.800 ;
        RECT 54.200 66.200 54.500 75.800 ;
        RECT 58.200 75.200 58.500 81.800 ;
        RECT 61.400 77.800 61.800 78.200 ;
        RECT 58.200 74.800 58.600 75.200 ;
        RECT 59.000 74.800 59.400 75.200 ;
        RECT 60.600 74.800 61.000 75.200 ;
        RECT 58.200 70.200 58.500 74.800 ;
        RECT 59.000 74.200 59.300 74.800 ;
        RECT 60.600 74.200 60.900 74.800 ;
        RECT 61.400 74.200 61.700 77.800 ;
        RECT 65.400 75.200 65.700 82.800 ;
        RECT 66.200 81.800 66.600 82.200 ;
        RECT 66.200 75.200 66.500 81.800 ;
        RECT 67.800 76.200 68.100 83.800 ;
        RECT 67.800 75.800 68.200 76.200 ;
        RECT 69.400 75.200 69.700 85.800 ;
        RECT 70.200 81.200 70.500 86.800 ;
        RECT 79.800 86.200 80.100 86.800 ;
        RECT 73.400 86.100 73.800 86.200 ;
        RECT 74.200 86.100 74.600 86.200 ;
        RECT 73.400 85.800 74.600 86.100 ;
        RECT 76.600 86.100 77.000 86.200 ;
        RECT 77.400 86.100 77.800 86.200 ;
        RECT 76.600 85.800 77.800 86.100 ;
        RECT 79.800 85.800 80.200 86.200 ;
        RECT 80.600 85.800 81.000 86.200 ;
        RECT 80.600 85.200 80.900 85.800 ;
        RECT 71.000 85.100 71.400 85.200 ;
        RECT 71.800 85.100 72.200 85.200 ;
        RECT 71.000 84.800 72.200 85.100 ;
        RECT 78.200 84.800 78.600 85.200 ;
        RECT 80.600 84.800 81.000 85.200 ;
        RECT 78.200 84.200 78.500 84.800 ;
        RECT 72.600 83.800 73.000 84.200 ;
        RECT 78.200 83.800 78.600 84.200 ;
        RECT 72.600 83.200 72.900 83.800 ;
        RECT 72.600 82.800 73.000 83.200 ;
        RECT 70.200 80.800 70.600 81.200 ;
        RECT 72.600 80.800 73.000 81.200 ;
        RECT 72.600 79.200 72.900 80.800 ;
        RECT 81.400 79.200 81.700 93.800 ;
        RECT 83.000 93.100 83.400 93.200 ;
        RECT 83.800 93.100 84.200 93.200 ;
        RECT 83.000 92.800 84.200 93.100 ;
        RECT 84.600 92.800 85.000 93.200 ;
        RECT 82.200 89.800 82.600 90.200 ;
        RECT 82.200 87.200 82.500 89.800 ;
        RECT 83.000 89.100 83.400 89.200 ;
        RECT 83.800 89.100 84.200 89.200 ;
        RECT 83.000 88.800 84.200 89.100 ;
        RECT 82.200 86.800 82.600 87.200 ;
        RECT 83.000 86.800 83.400 87.200 ;
        RECT 83.000 85.200 83.300 86.800 ;
        RECT 83.800 85.800 84.200 86.200 ;
        RECT 83.800 85.200 84.100 85.800 ;
        RECT 83.000 84.800 83.400 85.200 ;
        RECT 83.800 84.800 84.200 85.200 ;
        RECT 83.000 83.200 83.300 84.800 ;
        RECT 83.000 82.800 83.400 83.200 ;
        RECT 72.600 78.800 73.000 79.200 ;
        RECT 76.600 79.100 77.000 79.200 ;
        RECT 77.400 79.100 77.800 79.200 ;
        RECT 76.600 78.800 77.800 79.100 ;
        RECT 80.600 78.800 81.000 79.200 ;
        RECT 81.400 78.800 81.800 79.200 ;
        RECT 70.200 76.100 70.600 76.200 ;
        RECT 71.000 76.100 71.400 76.200 ;
        RECT 70.200 75.800 71.400 76.100 ;
        RECT 71.800 75.800 72.200 76.200 ;
        RECT 62.200 74.800 62.600 75.200 ;
        RECT 63.000 74.800 63.400 75.200 ;
        RECT 65.400 74.800 65.800 75.200 ;
        RECT 66.200 74.800 66.600 75.200 ;
        RECT 67.000 75.100 67.400 75.200 ;
        RECT 67.800 75.100 68.200 75.200 ;
        RECT 67.000 74.800 68.200 75.100 ;
        RECT 69.400 74.800 69.800 75.200 ;
        RECT 71.000 74.800 71.400 75.200 ;
        RECT 62.200 74.200 62.500 74.800 ;
        RECT 63.000 74.200 63.300 74.800 ;
        RECT 71.000 74.200 71.300 74.800 ;
        RECT 71.800 74.200 72.100 75.800 ;
        RECT 80.600 75.200 80.900 78.800 ;
        RECT 83.800 76.800 84.200 77.200 ;
        RECT 83.800 75.200 84.100 76.800 ;
        RECT 72.600 75.100 73.000 75.200 ;
        RECT 73.400 75.100 73.800 75.200 ;
        RECT 72.600 74.800 73.800 75.100 ;
        RECT 74.200 74.800 74.600 75.200 ;
        RECT 75.000 74.800 75.400 75.200 ;
        RECT 75.800 75.100 76.200 75.200 ;
        RECT 76.600 75.100 77.000 75.200 ;
        RECT 75.800 74.800 77.000 75.100 ;
        RECT 78.200 75.100 78.600 75.200 ;
        RECT 79.000 75.100 79.400 75.200 ;
        RECT 78.200 74.800 79.400 75.100 ;
        RECT 80.600 74.800 81.000 75.200 ;
        RECT 82.200 74.800 82.600 75.200 ;
        RECT 83.800 74.800 84.200 75.200 ;
        RECT 59.000 73.800 59.400 74.200 ;
        RECT 60.600 73.800 61.000 74.200 ;
        RECT 61.400 73.800 61.800 74.200 ;
        RECT 62.200 73.800 62.600 74.200 ;
        RECT 63.000 73.800 63.400 74.200 ;
        RECT 64.600 73.800 65.000 74.200 ;
        RECT 65.400 74.100 65.800 74.200 ;
        RECT 66.200 74.100 66.600 74.200 ;
        RECT 65.400 73.800 66.600 74.100 ;
        RECT 67.800 74.100 68.200 74.200 ;
        RECT 68.600 74.100 69.000 74.200 ;
        RECT 67.800 73.800 69.000 74.100 ;
        RECT 71.000 73.800 71.400 74.200 ;
        RECT 71.800 73.800 72.200 74.200 ;
        RECT 60.600 72.800 61.000 73.200 ;
        RECT 60.600 72.200 60.900 72.800 ;
        RECT 60.600 71.800 61.000 72.200 ;
        RECT 58.200 69.800 58.600 70.200 ;
        RECT 58.200 69.100 58.600 69.200 ;
        RECT 59.000 69.100 59.400 69.200 ;
        RECT 58.200 68.800 59.400 69.100 ;
        RECT 55.000 67.800 55.400 68.200 ;
        RECT 59.000 67.800 59.400 68.200 ;
        RECT 55.000 67.200 55.300 67.800 ;
        RECT 55.000 66.800 55.400 67.200 ;
        RECT 57.400 66.800 57.800 67.200 ;
        RECT 54.200 65.800 54.600 66.200 ;
        RECT 56.600 65.800 57.000 66.200 ;
        RECT 54.200 65.200 54.500 65.800 ;
        RECT 56.600 65.200 56.900 65.800 ;
        RECT 54.200 64.800 54.600 65.200 ;
        RECT 55.000 65.100 55.400 65.200 ;
        RECT 55.800 65.100 56.200 65.200 ;
        RECT 55.000 64.800 56.200 65.100 ;
        RECT 56.600 64.800 57.000 65.200 ;
        RECT 57.400 58.200 57.700 66.800 ;
        RECT 58.200 64.800 58.600 65.200 ;
        RECT 58.200 64.200 58.500 64.800 ;
        RECT 58.200 63.800 58.600 64.200 ;
        RECT 57.400 57.800 57.800 58.200 ;
        RECT 55.800 57.100 56.200 57.200 ;
        RECT 56.600 57.100 57.000 57.200 ;
        RECT 55.800 56.800 57.000 57.100 ;
        RECT 55.800 55.800 56.200 56.200 ;
        RECT 55.800 55.200 56.100 55.800 ;
        RECT 55.800 54.800 56.200 55.200 ;
        RECT 53.400 53.800 53.800 54.200 ;
        RECT 55.000 53.800 55.400 54.200 ;
        RECT 51.800 48.800 52.200 49.200 ;
        RECT 53.400 48.800 53.800 49.200 ;
        RECT 51.000 46.800 51.400 47.200 ;
        RECT 43.800 39.200 44.100 42.800 ;
        RECT 51.000 42.200 51.300 46.800 ;
        RECT 51.800 46.200 52.100 48.800 ;
        RECT 51.800 45.800 52.200 46.200 ;
        RECT 53.400 45.200 53.700 48.800 ;
        RECT 54.200 46.800 54.600 47.200 ;
        RECT 52.600 44.800 53.000 45.200 ;
        RECT 53.400 44.800 53.800 45.200 ;
        RECT 51.000 41.800 51.400 42.200 ;
        RECT 43.800 38.800 44.200 39.200 ;
        RECT 42.200 36.800 43.300 37.100 ;
        RECT 51.800 37.800 52.200 38.200 ;
        RECT 39.800 35.800 40.200 36.200 ;
        RECT 39.800 35.200 40.100 35.800 ;
        RECT 39.800 34.800 40.200 35.200 ;
        RECT 40.600 34.800 41.000 35.200 ;
        RECT 40.600 34.200 40.900 34.800 ;
        RECT 40.600 33.800 41.000 34.200 ;
        RECT 42.200 33.200 42.500 36.800 ;
        RECT 43.000 35.800 43.400 36.200 ;
        RECT 45.400 36.100 45.800 36.200 ;
        RECT 46.200 36.100 46.600 36.200 ;
        RECT 45.400 35.800 46.600 36.100 ;
        RECT 47.800 35.800 48.200 36.200 ;
        RECT 43.000 34.200 43.300 35.800 ;
        RECT 47.800 35.200 48.100 35.800 ;
        RECT 43.800 34.800 44.200 35.200 ;
        RECT 46.200 34.800 46.600 35.200 ;
        RECT 47.800 34.800 48.200 35.200 ;
        RECT 51.000 34.800 51.400 35.200 ;
        RECT 43.800 34.200 44.100 34.800 ;
        RECT 43.000 33.800 43.400 34.200 ;
        RECT 43.800 33.800 44.200 34.200 ;
        RECT 46.200 33.200 46.500 34.800 ;
        RECT 47.000 33.800 47.400 34.200 ;
        RECT 48.600 33.800 49.000 34.200 ;
        RECT 38.200 32.800 38.600 33.200 ;
        RECT 39.000 32.800 39.400 33.200 ;
        RECT 42.200 32.800 42.600 33.200 ;
        RECT 46.200 32.800 46.600 33.200 ;
        RECT 39.000 32.200 39.300 32.800 ;
        RECT 47.000 32.200 47.300 33.800 ;
        RECT 48.600 33.200 48.900 33.800 ;
        RECT 48.600 32.800 49.000 33.200 ;
        RECT 33.400 31.800 33.800 32.200 ;
        RECT 39.000 31.800 39.400 32.200 ;
        RECT 41.400 31.800 41.800 32.200 ;
        RECT 47.000 31.800 47.400 32.200 ;
        RECT 41.400 30.200 41.700 31.800 ;
        RECT 51.000 30.200 51.300 34.800 ;
        RECT 51.800 34.200 52.100 37.800 ;
        RECT 51.800 33.800 52.200 34.200 ;
        RECT 41.400 29.800 41.800 30.200 ;
        RECT 51.000 29.800 51.400 30.200 ;
        RECT 31.000 28.800 31.400 29.200 ;
        RECT 34.200 28.800 34.600 29.200 ;
        RECT 31.000 25.200 31.300 28.800 ;
        RECT 31.800 28.100 32.200 28.200 ;
        RECT 32.600 28.100 33.000 28.200 ;
        RECT 31.800 27.800 33.000 28.100 ;
        RECT 34.200 27.200 34.500 28.800 ;
        RECT 34.200 26.800 34.600 27.200 ;
        RECT 32.600 26.100 33.000 26.200 ;
        RECT 33.400 26.100 33.800 26.200 ;
        RECT 32.600 25.800 33.800 26.100 ;
        RECT 31.000 24.800 31.400 25.200 ;
        RECT 24.600 17.100 25.000 17.200 ;
        RECT 25.400 17.100 25.800 17.200 ;
        RECT 24.600 16.800 25.800 17.100 ;
        RECT 30.200 16.800 30.600 17.200 ;
        RECT 31.800 16.800 32.200 17.200 ;
        RECT 26.200 15.800 26.600 16.200 ;
        RECT 28.600 16.100 29.000 16.200 ;
        RECT 29.400 16.100 29.800 16.200 ;
        RECT 28.600 15.800 29.800 16.100 ;
        RECT 26.200 15.200 26.500 15.800 ;
        RECT 26.200 14.800 26.600 15.200 ;
        RECT 27.000 15.100 27.400 15.200 ;
        RECT 27.800 15.100 28.200 15.200 ;
        RECT 27.000 14.800 28.200 15.100 ;
        RECT 30.200 14.200 30.500 16.800 ;
        RECT 31.800 15.200 32.100 16.800 ;
        RECT 31.800 14.800 32.200 15.200 ;
        RECT 32.600 14.200 32.900 25.800 ;
        RECT 34.200 17.200 34.500 26.800 ;
        RECT 35.000 25.100 35.400 27.900 ;
        RECT 35.800 27.800 36.200 28.200 ;
        RECT 35.800 27.200 36.100 27.800 ;
        RECT 35.800 26.800 36.200 27.200 ;
        RECT 36.600 23.100 37.000 28.900 ;
        RECT 39.800 26.800 40.200 27.200 ;
        RECT 38.200 25.800 38.600 26.200 ;
        RECT 38.200 25.200 38.500 25.800 ;
        RECT 38.200 24.800 38.600 25.200 ;
        RECT 37.400 19.100 37.800 19.200 ;
        RECT 38.200 19.100 38.600 19.200 ;
        RECT 37.400 18.800 38.600 19.100 ;
        RECT 34.200 16.800 34.600 17.200 ;
        RECT 39.800 16.200 40.100 26.800 ;
        RECT 41.400 23.100 41.800 28.900 ;
        RECT 43.800 28.800 44.200 29.200 ;
        RECT 46.200 28.800 46.600 29.200 ;
        RECT 43.800 28.200 44.100 28.800 ;
        RECT 43.800 27.800 44.200 28.200 ;
        RECT 44.600 27.100 45.000 27.200 ;
        RECT 45.400 27.100 45.800 27.200 ;
        RECT 44.600 26.800 45.800 27.100 ;
        RECT 46.200 26.200 46.500 28.800 ;
        RECT 49.400 27.800 49.800 28.200 ;
        RECT 49.400 27.200 49.700 27.800 ;
        RECT 47.800 26.800 48.200 27.200 ;
        RECT 49.400 26.800 49.800 27.200 ;
        RECT 50.200 26.800 50.600 27.200 ;
        RECT 45.400 26.100 45.800 26.200 ;
        RECT 46.200 26.100 46.600 26.200 ;
        RECT 45.400 25.800 46.600 26.100 ;
        RECT 47.800 25.200 48.100 26.800 ;
        RECT 50.200 25.200 50.500 26.800 ;
        RECT 45.400 24.800 45.800 25.200 ;
        RECT 47.800 25.100 48.200 25.200 ;
        RECT 48.600 25.100 49.000 25.200 ;
        RECT 47.800 24.800 49.000 25.100 ;
        RECT 50.200 24.800 50.600 25.200 ;
        RECT 45.400 24.200 45.700 24.800 ;
        RECT 45.400 23.800 45.800 24.200 ;
        RECT 49.400 18.100 49.800 18.200 ;
        RECT 50.200 18.100 50.600 18.200 ;
        RECT 34.200 15.800 34.600 16.200 ;
        RECT 39.800 15.800 40.200 16.200 ;
        RECT 34.200 15.200 34.500 15.800 ;
        RECT 34.200 14.800 34.600 15.200 ;
        RECT 38.200 14.800 38.600 15.200 ;
        RECT 38.200 14.200 38.500 14.800 ;
        RECT 25.400 14.100 25.800 14.200 ;
        RECT 26.200 14.100 26.600 14.200 ;
        RECT 25.400 13.800 26.600 14.100 ;
        RECT 30.200 13.800 30.600 14.200 ;
        RECT 31.000 14.100 31.400 14.200 ;
        RECT 31.800 14.100 32.200 14.200 ;
        RECT 31.000 13.800 32.200 14.100 ;
        RECT 32.600 13.800 33.000 14.200 ;
        RECT 35.800 13.800 36.200 14.200 ;
        RECT 36.600 13.800 37.000 14.200 ;
        RECT 38.200 13.800 38.600 14.200 ;
        RECT 35.800 13.200 36.100 13.800 ;
        RECT 36.600 13.200 36.900 13.800 ;
        RECT 39.800 13.200 40.100 15.800 ;
        RECT 35.800 12.800 36.200 13.200 ;
        RECT 36.600 12.800 37.000 13.200 ;
        RECT 39.000 12.800 39.400 13.200 ;
        RECT 39.800 12.800 40.200 13.200 ;
        RECT 40.600 13.100 41.000 15.900 ;
        RECT 41.400 12.800 41.800 13.200 ;
        RECT 39.000 12.200 39.300 12.800 ;
        RECT 33.400 11.800 33.800 12.200 ;
        RECT 39.000 11.800 39.400 12.200 ;
        RECT 39.800 11.800 40.200 12.200 ;
        RECT 26.200 10.800 26.600 11.200 ;
        RECT 28.600 10.800 29.000 11.200 ;
        RECT 24.600 9.800 25.000 10.200 ;
        RECT 6.200 8.800 6.600 9.200 ;
        RECT 14.200 6.800 14.600 7.200 ;
        RECT 14.200 6.200 14.500 6.800 ;
        RECT 14.200 5.800 14.600 6.200 ;
        RECT 15.000 5.100 15.400 7.900 ;
        RECT 15.800 6.800 16.200 7.200 ;
        RECT 15.800 6.200 16.100 6.800 ;
        RECT 15.800 5.800 16.200 6.200 ;
        RECT 16.600 3.100 17.000 8.900 ;
        RECT 18.200 6.100 18.600 6.200 ;
        RECT 19.000 6.100 19.400 6.200 ;
        RECT 18.200 5.800 19.400 6.100 ;
        RECT 21.400 3.100 21.800 8.900 ;
        RECT 24.600 8.200 24.900 9.800 ;
        RECT 24.600 7.800 25.000 8.200 ;
        RECT 26.200 6.200 26.500 10.800 ;
        RECT 28.600 7.200 28.900 10.800 ;
        RECT 27.000 6.800 27.400 7.200 ;
        RECT 28.600 6.800 29.000 7.200 ;
        RECT 27.000 6.200 27.300 6.800 ;
        RECT 26.200 5.800 26.600 6.200 ;
        RECT 27.000 5.800 27.400 6.200 ;
        RECT 28.600 6.100 29.000 6.200 ;
        RECT 29.400 6.100 29.800 6.200 ;
        RECT 28.600 5.800 29.800 6.100 ;
        RECT 30.200 5.100 30.600 7.900 ;
        RECT 31.000 6.800 31.400 7.200 ;
        RECT 31.000 6.200 31.300 6.800 ;
        RECT 31.000 5.800 31.400 6.200 ;
        RECT 31.800 3.100 32.200 8.900 ;
        RECT 33.400 6.200 33.700 11.800 ;
        RECT 39.000 9.200 39.300 11.800 ;
        RECT 33.400 5.800 33.800 6.200 ;
        RECT 36.600 3.100 37.000 8.900 ;
        RECT 39.000 8.800 39.400 9.200 ;
        RECT 39.800 5.200 40.100 11.800 ;
        RECT 41.400 10.100 41.700 12.800 ;
        RECT 42.200 12.100 42.600 17.900 ;
        RECT 43.800 15.100 44.200 15.200 ;
        RECT 44.600 15.100 45.000 15.200 ;
        RECT 43.800 14.800 45.000 15.100 ;
        RECT 43.000 13.800 43.400 14.200 ;
        RECT 43.800 13.800 44.200 14.200 ;
        RECT 41.400 9.800 42.500 10.100 ;
        RECT 41.400 8.800 41.800 9.200 ;
        RECT 41.400 6.200 41.700 8.800 ;
        RECT 42.200 7.200 42.500 9.800 ;
        RECT 43.000 9.200 43.300 13.800 ;
        RECT 43.000 8.800 43.400 9.200 ;
        RECT 42.200 6.800 42.600 7.200 ;
        RECT 43.800 6.200 44.100 13.800 ;
        RECT 47.000 12.100 47.400 17.900 ;
        RECT 49.400 17.800 50.600 18.100 ;
        RECT 51.800 16.800 52.200 17.200 ;
        RECT 51.800 14.200 52.100 16.800 ;
        RECT 52.600 15.200 52.900 44.800 ;
        RECT 53.400 43.800 53.800 44.200 ;
        RECT 54.200 44.100 54.500 46.800 ;
        RECT 55.000 45.200 55.300 53.800 ;
        RECT 56.600 52.800 57.000 53.200 ;
        RECT 56.600 49.200 56.900 52.800 ;
        RECT 57.400 51.200 57.700 57.800 ;
        RECT 58.200 56.800 58.600 57.200 ;
        RECT 58.200 56.200 58.500 56.800 ;
        RECT 58.200 55.800 58.600 56.200 ;
        RECT 59.000 55.100 59.300 67.800 ;
        RECT 59.800 66.800 60.200 67.200 ;
        RECT 59.800 61.200 60.100 66.800 ;
        RECT 60.600 65.100 61.000 67.900 ;
        RECT 61.400 66.800 61.800 67.200 ;
        RECT 59.800 60.800 60.200 61.200 ;
        RECT 60.600 58.800 61.000 59.200 ;
        RECT 60.600 56.200 60.900 58.800 ;
        RECT 60.600 55.800 61.000 56.200 ;
        RECT 58.200 54.800 59.300 55.100 ;
        RECT 59.800 54.800 60.200 55.200 ;
        RECT 57.400 50.800 57.800 51.200 ;
        RECT 56.600 48.800 57.000 49.200 ;
        RECT 57.400 45.800 57.800 46.200 ;
        RECT 55.000 44.800 55.400 45.200 ;
        RECT 56.600 44.800 57.000 45.200 ;
        RECT 54.200 43.800 55.300 44.100 ;
        RECT 53.400 39.200 53.700 43.800 ;
        RECT 55.000 39.200 55.300 43.800 ;
        RECT 56.600 43.200 56.900 44.800 ;
        RECT 56.600 42.800 57.000 43.200 ;
        RECT 57.400 40.200 57.700 45.800 ;
        RECT 57.400 39.800 57.800 40.200 ;
        RECT 58.200 39.200 58.500 54.800 ;
        RECT 59.800 54.200 60.100 54.800 ;
        RECT 59.800 53.800 60.200 54.200 ;
        RECT 59.000 50.800 59.400 51.200 ;
        RECT 59.000 49.200 59.300 50.800 ;
        RECT 60.600 49.200 60.900 55.800 ;
        RECT 59.000 48.800 59.400 49.200 ;
        RECT 60.600 48.800 61.000 49.200 ;
        RECT 60.600 45.100 61.000 47.900 ;
        RECT 61.400 47.200 61.700 66.800 ;
        RECT 62.200 63.100 62.600 68.900 ;
        RECT 64.600 68.200 64.900 73.800 ;
        RECT 67.800 73.100 68.200 73.200 ;
        RECT 68.600 73.100 69.000 73.200 ;
        RECT 67.800 72.800 69.000 73.100 ;
        RECT 65.400 68.800 65.800 69.200 ;
        RECT 71.000 69.100 71.400 69.200 ;
        RECT 71.800 69.100 72.200 69.200 ;
        RECT 64.600 67.800 65.000 68.200 ;
        RECT 65.400 66.200 65.700 68.800 ;
        RECT 65.400 65.800 65.800 66.200 ;
        RECT 67.000 63.100 67.400 68.900 ;
        RECT 71.000 68.800 72.200 69.100 ;
        RECT 69.400 68.100 69.800 68.200 ;
        RECT 70.200 68.100 70.600 68.200 ;
        RECT 69.400 67.800 70.600 68.100 ;
        RECT 72.600 68.100 73.000 68.200 ;
        RECT 73.400 68.100 73.800 68.200 ;
        RECT 72.600 67.800 73.800 68.100 ;
        RECT 70.200 67.100 70.600 67.200 ;
        RECT 71.000 67.100 71.400 67.200 ;
        RECT 70.200 66.800 71.400 67.100 ;
        RECT 70.200 66.100 70.600 66.200 ;
        RECT 71.000 66.100 71.400 66.200 ;
        RECT 70.200 65.800 71.400 66.100 ;
        RECT 73.400 65.200 73.700 67.800 ;
        RECT 73.400 64.800 73.800 65.200 ;
        RECT 74.200 63.200 74.500 74.800 ;
        RECT 75.000 74.200 75.300 74.800 ;
        RECT 82.200 74.200 82.500 74.800 ;
        RECT 75.000 73.800 75.400 74.200 ;
        RECT 75.800 73.800 76.200 74.200 ;
        RECT 78.200 74.100 78.600 74.200 ;
        RECT 79.000 74.100 79.400 74.200 ;
        RECT 78.200 73.800 79.400 74.100 ;
        RECT 79.800 73.800 80.200 74.200 ;
        RECT 82.200 73.800 82.600 74.200 ;
        RECT 83.000 73.800 83.400 74.200 ;
        RECT 83.800 73.800 84.200 74.200 ;
        RECT 75.800 73.200 76.100 73.800 ;
        RECT 79.800 73.200 80.100 73.800 ;
        RECT 83.000 73.200 83.300 73.800 ;
        RECT 75.800 72.800 76.200 73.200 ;
        RECT 79.800 72.800 80.200 73.200 ;
        RECT 80.600 72.800 81.000 73.200 ;
        RECT 83.000 72.800 83.400 73.200 ;
        RECT 79.000 69.800 79.400 70.200 ;
        RECT 79.000 69.200 79.300 69.800 ;
        RECT 75.800 68.800 76.200 69.200 ;
        RECT 79.000 68.800 79.400 69.200 ;
        RECT 75.000 66.800 75.400 67.200 ;
        RECT 75.000 66.200 75.300 66.800 ;
        RECT 75.800 66.200 76.100 68.800 ;
        RECT 75.000 65.800 75.400 66.200 ;
        RECT 75.800 65.800 76.200 66.200 ;
        RECT 74.200 62.800 74.600 63.200 ;
        RECT 66.200 61.800 66.600 62.200 ;
        RECT 62.200 60.800 62.600 61.200 ;
        RECT 62.200 59.200 62.500 60.800 ;
        RECT 62.200 58.800 62.600 59.200 ;
        RECT 63.000 57.800 63.400 58.200 ;
        RECT 63.000 57.200 63.300 57.800 ;
        RECT 63.000 56.800 63.400 57.200 ;
        RECT 63.000 55.200 63.300 56.800 ;
        RECT 62.200 54.800 62.600 55.200 ;
        RECT 63.000 54.800 63.400 55.200 ;
        RECT 65.400 54.800 65.800 55.200 ;
        RECT 62.200 54.200 62.500 54.800 ;
        RECT 65.400 54.200 65.700 54.800 ;
        RECT 62.200 53.800 62.600 54.200 ;
        RECT 63.000 54.100 63.400 54.200 ;
        RECT 63.800 54.100 64.200 54.200 ;
        RECT 63.000 53.800 64.200 54.100 ;
        RECT 64.600 53.800 65.000 54.200 ;
        RECT 65.400 53.800 65.800 54.200 ;
        RECT 61.400 46.800 61.800 47.200 ;
        RECT 61.400 46.200 61.700 46.800 ;
        RECT 61.400 45.800 61.800 46.200 ;
        RECT 62.200 43.100 62.600 48.900 ;
        RECT 64.600 48.200 64.900 53.800 ;
        RECT 66.200 53.200 66.500 61.800 ;
        RECT 66.200 52.800 66.600 53.200 ;
        RECT 67.000 53.100 67.400 55.900 ;
        RECT 68.600 52.100 69.000 57.900 ;
        RECT 70.200 55.100 70.600 55.200 ;
        RECT 71.000 55.100 71.400 55.200 ;
        RECT 70.200 54.800 71.400 55.100 ;
        RECT 71.000 53.800 71.400 54.200 ;
        RECT 64.600 47.800 65.000 48.200 ;
        RECT 65.400 45.800 65.800 46.200 ;
        RECT 53.400 38.800 53.800 39.200 ;
        RECT 55.000 38.800 55.400 39.200 ;
        RECT 58.200 38.800 58.600 39.200 ;
        RECT 61.400 37.800 61.800 38.200 ;
        RECT 55.800 35.800 56.200 36.200 ;
        RECT 59.000 36.100 59.400 36.200 ;
        RECT 59.800 36.100 60.200 36.200 ;
        RECT 59.000 35.800 60.200 36.100 ;
        RECT 55.800 35.200 56.100 35.800 ;
        RECT 61.400 35.200 61.700 37.800 ;
        RECT 65.400 36.200 65.700 45.800 ;
        RECT 67.000 43.100 67.400 48.900 ;
        RECT 70.200 45.100 70.600 47.900 ;
        RECT 71.000 47.200 71.300 53.800 ;
        RECT 73.400 52.100 73.800 57.900 ;
        RECT 75.000 54.200 75.300 65.800 ;
        RECT 79.000 64.800 79.400 65.200 ;
        RECT 77.400 63.800 77.800 64.200 ;
        RECT 77.400 63.200 77.700 63.800 ;
        RECT 77.400 62.800 77.800 63.200 ;
        RECT 79.000 60.200 79.300 64.800 ;
        RECT 79.000 59.800 79.400 60.200 ;
        RECT 75.800 58.100 76.200 58.200 ;
        RECT 76.600 58.100 77.000 58.200 ;
        RECT 75.800 57.800 77.000 58.100 ;
        RECT 77.400 56.100 77.800 56.200 ;
        RECT 76.600 55.800 77.800 56.100 ;
        RECT 79.800 55.800 80.200 56.200 ;
        RECT 76.600 55.200 76.900 55.800 ;
        RECT 79.800 55.200 80.100 55.800 ;
        RECT 76.600 54.800 77.000 55.200 ;
        RECT 77.400 54.800 77.800 55.200 ;
        RECT 79.800 54.800 80.200 55.200 ;
        RECT 75.000 53.800 75.400 54.200 ;
        RECT 76.600 53.800 77.000 54.200 ;
        RECT 76.600 53.200 76.900 53.800 ;
        RECT 76.600 52.800 77.000 53.200 ;
        RECT 71.000 46.800 71.400 47.200 ;
        RECT 71.000 46.200 71.300 46.800 ;
        RECT 71.000 45.800 71.400 46.200 ;
        RECT 69.400 42.800 69.800 43.200 ;
        RECT 71.800 43.100 72.200 48.900 ;
        RECT 75.000 47.800 75.400 48.200 ;
        RECT 75.000 46.200 75.300 47.800 ;
        RECT 75.000 45.800 75.400 46.200 ;
        RECT 75.000 43.800 75.400 44.200 ;
        RECT 69.400 42.200 69.700 42.800 ;
        RECT 69.400 41.800 69.800 42.200 ;
        RECT 68.600 38.800 69.000 39.200 ;
        RECT 68.600 36.200 68.900 38.800 ;
        RECT 63.000 36.100 63.400 36.200 ;
        RECT 63.800 36.100 64.200 36.200 ;
        RECT 63.000 35.800 64.200 36.100 ;
        RECT 64.600 35.800 65.000 36.200 ;
        RECT 65.400 35.800 65.800 36.200 ;
        RECT 67.000 35.800 67.400 36.200 ;
        RECT 68.600 35.800 69.000 36.200 ;
        RECT 64.600 35.200 64.900 35.800 ;
        RECT 67.000 35.200 67.300 35.800 ;
        RECT 55.800 34.800 56.200 35.200 ;
        RECT 61.400 34.800 61.800 35.200 ;
        RECT 64.600 34.800 65.000 35.200 ;
        RECT 65.400 35.100 65.800 35.200 ;
        RECT 66.200 35.100 66.600 35.200 ;
        RECT 65.400 34.800 66.600 35.100 ;
        RECT 67.000 34.800 67.400 35.200 ;
        RECT 68.600 34.200 68.900 35.800 ;
        RECT 53.400 33.800 53.800 34.200 ;
        RECT 58.200 33.800 58.600 34.200 ;
        RECT 61.400 33.800 61.800 34.200 ;
        RECT 62.200 33.800 62.600 34.200 ;
        RECT 65.400 34.100 65.800 34.200 ;
        RECT 66.200 34.100 66.600 34.200 ;
        RECT 65.400 33.800 66.600 34.100 ;
        RECT 68.600 33.800 69.000 34.200 ;
        RECT 69.400 34.100 69.700 41.800 ;
        RECT 75.000 41.200 75.300 43.800 ;
        RECT 76.600 43.100 77.000 48.900 ;
        RECT 77.400 47.200 77.700 54.800 ;
        RECT 80.600 54.100 80.900 72.800 ;
        RECT 83.800 72.100 84.100 73.800 ;
        RECT 83.000 71.800 84.100 72.100 ;
        RECT 81.400 65.800 81.800 66.200 ;
        RECT 81.400 65.200 81.700 65.800 ;
        RECT 81.400 64.800 81.800 65.200 ;
        RECT 79.800 53.800 80.900 54.100 ;
        RECT 81.400 57.800 81.800 58.200 ;
        RECT 81.400 54.200 81.700 57.800 ;
        RECT 83.000 57.200 83.300 71.800 ;
        RECT 84.600 69.200 84.900 92.800 ;
        RECT 85.400 91.200 85.700 93.800 ;
        RECT 85.400 90.800 85.800 91.200 ;
        RECT 87.000 90.200 87.300 94.800 ;
        RECT 91.800 94.200 92.100 97.800 ;
        RECT 93.400 96.200 93.700 98.800 ;
        RECT 93.400 95.800 93.800 96.200 ;
        RECT 92.600 95.100 93.000 95.200 ;
        RECT 93.400 95.100 93.800 95.200 ;
        RECT 92.600 94.800 93.800 95.100 ;
        RECT 90.200 94.100 90.600 94.200 ;
        RECT 90.200 93.800 91.300 94.100 ;
        RECT 91.800 93.800 92.200 94.200 ;
        RECT 91.000 93.200 91.300 93.800 ;
        RECT 89.400 93.100 89.800 93.200 ;
        RECT 90.200 93.100 90.600 93.200 ;
        RECT 89.400 92.800 90.600 93.100 ;
        RECT 91.000 92.800 91.400 93.200 ;
        RECT 88.600 91.800 89.000 92.200 ;
        RECT 93.400 91.800 93.800 92.200 ;
        RECT 88.600 91.200 88.900 91.800 ;
        RECT 88.600 90.800 89.000 91.200 ;
        RECT 87.000 89.800 87.400 90.200 ;
        RECT 85.400 88.800 85.800 89.200 ;
        RECT 89.400 89.100 89.800 89.200 ;
        RECT 90.200 89.100 90.600 89.200 ;
        RECT 89.400 88.800 90.600 89.100 ;
        RECT 85.400 86.200 85.700 88.800 ;
        RECT 93.400 88.200 93.700 91.800 ;
        RECT 93.400 87.800 93.800 88.200 ;
        RECT 86.200 86.800 86.600 87.200 ;
        RECT 87.000 87.100 87.400 87.200 ;
        RECT 87.800 87.100 88.200 87.200 ;
        RECT 87.000 86.800 88.200 87.100 ;
        RECT 91.800 87.100 92.200 87.200 ;
        RECT 92.600 87.100 93.000 87.200 ;
        RECT 91.800 86.800 93.000 87.100 ;
        RECT 85.400 85.800 85.800 86.200 ;
        RECT 86.200 84.200 86.500 86.800 ;
        RECT 87.000 85.800 87.400 86.200 ;
        RECT 91.000 85.800 91.400 86.200 ;
        RECT 86.200 83.800 86.600 84.200 ;
        RECT 86.200 77.800 86.600 78.200 ;
        RECT 86.200 76.200 86.500 77.800 ;
        RECT 86.200 75.800 86.600 76.200 ;
        RECT 85.400 71.800 85.800 72.200 ;
        RECT 84.600 68.800 85.000 69.200 ;
        RECT 83.800 67.100 84.200 67.200 ;
        RECT 84.600 67.100 85.000 67.200 ;
        RECT 83.800 66.800 85.000 67.100 ;
        RECT 84.600 66.100 85.000 66.200 ;
        RECT 85.400 66.100 85.700 71.800 ;
        RECT 87.000 69.200 87.300 85.800 ;
        RECT 91.000 84.200 91.300 85.800 ;
        RECT 94.200 85.200 94.500 101.800 ;
        RECT 96.600 96.100 96.900 101.800 ;
        RECT 97.400 99.200 97.700 104.800 ;
        RECT 98.200 104.200 98.500 106.800 ;
        RECT 99.800 105.200 100.100 106.800 ;
        RECT 99.800 104.800 100.200 105.200 ;
        RECT 98.200 103.800 98.600 104.200 ;
        RECT 97.400 98.800 97.800 99.200 ;
        RECT 95.800 95.800 96.900 96.100 ;
        RECT 95.800 95.200 96.100 95.800 ;
        RECT 95.800 94.800 96.200 95.200 ;
        RECT 96.600 94.800 97.000 95.200 ;
        RECT 96.600 94.200 96.900 94.800 ;
        RECT 96.600 93.800 97.000 94.200 ;
        RECT 96.600 87.200 96.900 93.800 ;
        RECT 97.400 91.800 97.800 92.200 ;
        RECT 96.600 86.800 97.000 87.200 ;
        RECT 94.200 84.800 94.600 85.200 ;
        RECT 91.000 83.800 91.400 84.200 ;
        RECT 94.200 82.200 94.500 84.800 ;
        RECT 96.600 84.200 96.900 86.800 ;
        RECT 96.600 83.800 97.000 84.200 ;
        RECT 91.800 81.800 92.200 82.200 ;
        RECT 93.400 81.800 93.800 82.200 ;
        RECT 94.200 81.800 94.600 82.200 ;
        RECT 95.800 81.800 96.200 82.200 ;
        RECT 91.800 79.200 92.100 81.800 ;
        RECT 91.800 78.800 92.200 79.200 ;
        RECT 93.400 77.200 93.700 81.800 ;
        RECT 94.200 80.800 94.600 81.200 ;
        RECT 91.800 76.800 92.200 77.200 ;
        RECT 93.400 76.800 93.800 77.200 ;
        RECT 87.800 75.800 88.200 76.200 ;
        RECT 88.600 75.800 89.000 76.200 ;
        RECT 87.800 73.100 88.100 75.800 ;
        RECT 88.600 74.200 88.900 75.800 ;
        RECT 89.400 74.800 89.800 75.200 ;
        RECT 91.000 74.800 91.400 75.200 ;
        RECT 89.400 74.200 89.700 74.800 ;
        RECT 91.000 74.200 91.300 74.800 ;
        RECT 88.600 73.800 89.000 74.200 ;
        RECT 89.400 73.800 89.800 74.200 ;
        RECT 90.200 73.800 90.600 74.200 ;
        RECT 91.000 73.800 91.400 74.200 ;
        RECT 90.200 73.100 90.500 73.800 ;
        RECT 87.800 72.800 90.500 73.100 ;
        RECT 87.800 72.100 88.200 72.200 ;
        RECT 88.600 72.100 89.000 72.200 ;
        RECT 87.800 71.800 89.000 72.100 ;
        RECT 90.200 71.800 90.600 72.200 ;
        RECT 87.800 70.800 88.200 71.200 ;
        RECT 87.800 69.200 88.100 70.800 ;
        RECT 87.000 68.800 87.400 69.200 ;
        RECT 87.800 68.800 88.200 69.200 ;
        RECT 87.000 67.800 87.400 68.200 ;
        RECT 87.000 67.200 87.300 67.800 ;
        RECT 87.000 66.800 87.400 67.200 ;
        RECT 90.200 66.200 90.500 71.800 ;
        RECT 91.800 66.200 92.100 76.800 ;
        RECT 92.600 75.100 93.000 75.200 ;
        RECT 93.400 75.100 93.800 75.200 ;
        RECT 92.600 74.800 93.800 75.100 ;
        RECT 93.400 73.800 93.800 74.200 ;
        RECT 93.400 69.200 93.700 73.800 ;
        RECT 94.200 73.200 94.500 80.800 ;
        RECT 95.800 77.200 96.100 81.800 ;
        RECT 97.400 80.200 97.700 91.800 ;
        RECT 98.200 88.200 98.500 103.800 ;
        RECT 99.000 97.800 99.400 98.200 ;
        RECT 99.000 95.200 99.300 97.800 ;
        RECT 99.000 94.800 99.400 95.200 ;
        RECT 99.000 94.200 99.300 94.800 ;
        RECT 99.000 93.800 99.400 94.200 ;
        RECT 99.800 93.800 100.200 94.200 ;
        RECT 98.200 87.800 98.600 88.200 ;
        RECT 99.000 86.800 99.400 87.200 ;
        RECT 99.000 86.200 99.300 86.800 ;
        RECT 99.000 85.800 99.400 86.200 ;
        RECT 97.400 79.800 97.800 80.200 ;
        RECT 99.800 78.200 100.100 93.800 ;
        RECT 100.600 88.200 100.900 124.800 ;
        RECT 102.200 113.800 102.600 114.200 ;
        RECT 102.200 113.200 102.500 113.800 ;
        RECT 102.200 112.800 102.600 113.200 ;
        RECT 102.200 112.200 102.500 112.800 ;
        RECT 102.200 111.800 102.600 112.200 ;
        RECT 103.800 106.200 104.100 137.800 ;
        RECT 105.400 135.200 105.700 137.800 ;
        RECT 105.400 134.800 105.800 135.200 ;
        RECT 106.200 134.800 106.600 135.200 ;
        RECT 108.600 135.100 109.000 135.200 ;
        RECT 109.400 135.100 109.800 135.200 ;
        RECT 108.600 134.800 109.800 135.100 ;
        RECT 104.600 133.800 105.000 134.200 ;
        RECT 104.600 131.200 104.900 133.800 ;
        RECT 104.600 130.800 105.000 131.200 ;
        RECT 104.600 127.100 105.000 127.200 ;
        RECT 105.400 127.100 105.800 127.200 ;
        RECT 104.600 126.800 105.800 127.100 ;
        RECT 104.600 126.100 105.000 126.200 ;
        RECT 105.400 126.100 105.800 126.200 ;
        RECT 104.600 125.800 105.800 126.100 ;
        RECT 106.200 125.200 106.500 134.800 ;
        RECT 110.200 134.200 110.500 143.800 ;
        RECT 115.800 140.200 116.100 143.800 ;
        RECT 118.200 143.200 118.500 145.800 ;
        RECT 119.000 144.200 119.300 147.800 ;
        RECT 121.400 146.100 121.800 146.200 ;
        RECT 122.200 146.100 122.600 146.200 ;
        RECT 121.400 145.800 122.600 146.100 ;
        RECT 123.800 145.200 124.100 150.800 ;
        RECT 124.600 150.200 124.900 155.800 ;
        RECT 125.400 151.800 125.800 152.200 ;
        RECT 124.600 149.800 125.000 150.200 ;
        RECT 125.400 149.200 125.700 151.800 ;
        RECT 125.400 148.800 125.800 149.200 ;
        RECT 124.600 145.800 125.000 146.200 ;
        RECT 120.600 144.800 121.000 145.200 ;
        RECT 123.800 144.800 124.200 145.200 ;
        RECT 120.600 144.200 120.900 144.800 ;
        RECT 119.000 143.800 119.400 144.200 ;
        RECT 120.600 143.800 121.000 144.200 ;
        RECT 122.200 144.100 122.600 144.200 ;
        RECT 123.000 144.100 123.400 144.200 ;
        RECT 122.200 143.800 123.400 144.100 ;
        RECT 124.600 143.200 124.900 145.800 ;
        RECT 125.400 145.200 125.700 148.800 ;
        RECT 127.000 146.200 127.300 171.800 ;
        RECT 128.600 167.200 128.900 171.800 ;
        RECT 140.600 170.200 140.900 173.800 ;
        RECT 141.400 172.100 141.800 177.900 ;
        RECT 142.200 172.100 142.600 178.900 ;
        RECT 143.000 172.100 143.400 178.900 ;
        RECT 146.200 174.800 146.600 175.200 ;
        RECT 151.000 174.800 151.400 175.200 ;
        RECT 146.200 174.200 146.500 174.800 ;
        RECT 151.000 174.200 151.300 174.800 ;
        RECT 146.200 173.800 146.600 174.200 ;
        RECT 148.600 173.800 149.000 174.200 ;
        RECT 151.000 173.800 151.400 174.200 ;
        RECT 143.800 172.800 144.200 173.200 ;
        RECT 140.600 169.800 141.000 170.200 ;
        RECT 130.100 167.500 130.500 167.900 ;
        RECT 131.000 167.500 133.100 167.800 ;
        RECT 133.400 167.500 133.800 167.900 ;
        RECT 128.600 166.800 129.000 167.200 ;
        RECT 129.400 166.800 129.800 167.200 ;
        RECT 128.600 165.800 129.000 166.200 ;
        RECT 127.800 157.800 128.200 158.200 ;
        RECT 127.800 146.200 128.100 157.800 ;
        RECT 128.600 151.200 128.900 165.800 ;
        RECT 129.400 156.200 129.700 166.800 ;
        RECT 130.100 165.100 130.400 167.500 ;
        RECT 131.000 167.400 131.400 167.500 ;
        RECT 132.700 167.400 133.100 167.500 ;
        RECT 133.500 167.100 133.800 167.500 ;
        RECT 131.400 166.800 133.800 167.100 ;
        RECT 134.200 167.800 134.600 168.200 ;
        RECT 134.200 167.200 134.500 167.800 ;
        RECT 134.200 166.800 134.600 167.200 ;
        RECT 131.400 166.700 131.800 166.800 ;
        RECT 133.500 165.100 133.800 166.800 ;
        RECT 130.100 164.700 130.500 165.100 ;
        RECT 133.400 164.700 133.800 165.100 ;
        RECT 131.800 164.100 132.200 164.200 ;
        RECT 132.600 164.100 133.000 164.200 ;
        RECT 131.800 163.800 133.000 164.100 ;
        RECT 140.600 162.100 141.000 168.900 ;
        RECT 141.400 162.100 141.800 168.900 ;
        RECT 142.200 162.100 142.600 168.900 ;
        RECT 143.000 163.100 143.400 168.900 ;
        RECT 143.800 168.200 144.100 172.800 ;
        RECT 143.800 167.800 144.200 168.200 ;
        RECT 144.600 163.100 145.000 168.900 ;
        RECT 145.400 166.800 145.800 167.200 ;
        RECT 145.400 164.200 145.700 166.800 ;
        RECT 145.400 163.800 145.800 164.200 ;
        RECT 146.200 163.100 146.600 168.900 ;
        RECT 147.000 162.100 147.400 168.900 ;
        RECT 147.800 162.100 148.200 168.900 ;
        RECT 148.600 166.200 148.900 173.800 ;
        RECT 151.000 172.800 151.400 173.200 ;
        RECT 148.600 165.800 149.000 166.200 ;
        RECT 129.400 155.800 129.800 156.200 ;
        RECT 128.600 150.800 129.000 151.200 ;
        RECT 129.400 146.200 129.700 155.800 ;
        RECT 130.200 152.100 130.600 158.900 ;
        RECT 131.000 152.100 131.400 158.900 ;
        RECT 131.800 152.100 132.200 158.900 ;
        RECT 132.600 152.100 133.000 157.900 ;
        RECT 133.400 153.800 133.800 154.200 ;
        RECT 133.400 153.200 133.700 153.800 ;
        RECT 133.400 152.800 133.800 153.200 ;
        RECT 134.200 152.100 134.600 157.900 ;
        RECT 135.000 153.800 135.400 154.200 ;
        RECT 133.400 150.800 133.800 151.200 ;
        RECT 133.400 149.200 133.700 150.800 ;
        RECT 135.000 150.200 135.300 153.800 ;
        RECT 135.800 152.100 136.200 157.900 ;
        RECT 136.600 152.100 137.000 158.900 ;
        RECT 137.400 152.100 137.800 158.900 ;
        RECT 138.200 154.800 138.600 155.200 ;
        RECT 147.000 154.800 147.400 155.200 ;
        RECT 138.200 153.200 138.500 154.800 ;
        RECT 147.000 153.200 147.300 154.800 ;
        RECT 138.200 152.800 138.600 153.200 ;
        RECT 147.000 152.800 147.400 153.200 ;
        RECT 143.000 152.100 143.400 152.200 ;
        RECT 143.800 152.100 144.200 152.200 ;
        RECT 143.000 151.800 144.200 152.100 ;
        RECT 146.200 151.800 146.600 152.200 ;
        RECT 147.800 152.100 148.200 158.900 ;
        RECT 148.600 152.100 149.000 158.900 ;
        RECT 149.400 152.100 149.800 158.900 ;
        RECT 150.200 152.100 150.600 157.900 ;
        RECT 151.000 154.200 151.300 172.800 ;
        RECT 153.400 172.100 153.800 178.900 ;
        RECT 154.200 172.100 154.600 178.900 ;
        RECT 155.000 172.100 155.400 177.900 ;
        RECT 155.800 173.800 156.200 174.200 ;
        RECT 155.800 169.100 156.100 173.800 ;
        RECT 156.600 172.100 157.000 177.900 ;
        RECT 157.400 173.800 157.800 174.200 ;
        RECT 157.400 173.200 157.700 173.800 ;
        RECT 157.400 172.800 157.800 173.200 ;
        RECT 158.200 172.100 158.600 177.900 ;
        RECT 159.000 172.100 159.400 178.900 ;
        RECT 159.800 172.100 160.200 178.900 ;
        RECT 160.600 172.100 161.000 178.900 ;
        RECT 161.400 174.800 161.800 175.200 ;
        RECT 177.400 174.800 177.800 175.200 ;
        RECT 161.400 169.200 161.700 174.800 ;
        RECT 173.400 173.800 173.800 174.200 ;
        RECT 173.400 173.200 173.700 173.800 ;
        RECT 173.400 172.800 173.800 173.200 ;
        RECT 165.400 171.800 165.800 172.200 ;
        RECT 156.600 169.100 157.000 169.200 ;
        RECT 155.800 168.800 157.000 169.100 ;
        RECT 161.400 168.800 161.800 169.200 ;
        RECT 155.000 167.500 155.400 167.900 ;
        RECT 155.700 167.500 157.800 167.800 ;
        RECT 158.300 167.500 158.700 167.900 ;
        RECT 154.200 166.800 154.600 167.200 ;
        RECT 155.000 167.100 155.300 167.500 ;
        RECT 155.700 167.400 156.100 167.500 ;
        RECT 157.400 167.400 157.800 167.500 ;
        RECT 155.000 166.800 157.400 167.100 ;
        RECT 154.200 166.200 154.500 166.800 ;
        RECT 154.200 165.800 154.600 166.200 ;
        RECT 155.000 165.100 155.300 166.800 ;
        RECT 157.000 166.700 157.400 166.800 ;
        RECT 158.400 165.100 158.700 167.500 ;
        RECT 160.500 167.500 160.900 167.900 ;
        RECT 161.400 167.500 163.500 167.800 ;
        RECT 163.800 167.500 164.200 167.900 ;
        RECT 159.000 166.800 159.400 167.200 ;
        RECT 159.800 166.800 160.200 167.200 ;
        RECT 159.000 166.200 159.300 166.800 ;
        RECT 159.000 165.800 159.400 166.200 ;
        RECT 155.000 164.700 155.400 165.100 ;
        RECT 158.300 164.700 158.700 165.100 ;
        RECT 151.000 153.800 151.400 154.200 ;
        RECT 151.000 153.200 151.300 153.800 ;
        RECT 151.000 152.800 151.400 153.200 ;
        RECT 151.800 152.100 152.200 157.900 ;
        RECT 152.600 153.800 153.000 154.200 ;
        RECT 135.800 150.800 136.200 151.200 ;
        RECT 135.000 149.800 135.400 150.200 ;
        RECT 133.400 148.800 133.800 149.200 ;
        RECT 135.800 148.200 136.100 150.800 ;
        RECT 140.600 149.800 141.000 150.200 ;
        RECT 140.600 149.200 140.900 149.800 ;
        RECT 140.600 148.800 141.000 149.200 ;
        RECT 143.000 148.800 143.400 149.200 ;
        RECT 130.200 148.100 130.600 148.200 ;
        RECT 131.000 148.100 131.400 148.200 ;
        RECT 130.200 147.800 131.400 148.100 ;
        RECT 135.800 147.800 136.200 148.200 ;
        RECT 139.000 147.500 139.400 147.900 ;
        RECT 139.700 147.500 141.800 147.800 ;
        RECT 142.300 147.500 142.700 147.900 ;
        RECT 136.600 147.100 137.000 147.200 ;
        RECT 137.400 147.100 137.800 147.200 ;
        RECT 136.600 146.800 137.800 147.100 ;
        RECT 138.200 146.800 138.600 147.200 ;
        RECT 139.000 147.100 139.300 147.500 ;
        RECT 139.700 147.400 140.100 147.500 ;
        RECT 141.400 147.400 141.800 147.500 ;
        RECT 139.000 146.800 141.400 147.100 ;
        RECT 127.000 145.800 127.400 146.200 ;
        RECT 127.800 145.800 128.200 146.200 ;
        RECT 129.400 145.800 129.800 146.200 ;
        RECT 131.800 145.800 132.200 146.200 ;
        RECT 135.000 145.800 135.400 146.200 ;
        RECT 136.600 146.100 137.000 146.200 ;
        RECT 137.400 146.100 137.800 146.200 ;
        RECT 136.600 145.800 137.800 146.100 ;
        RECT 127.000 145.200 127.300 145.800 ;
        RECT 127.800 145.200 128.100 145.800 ;
        RECT 125.400 144.800 125.800 145.200 ;
        RECT 127.000 144.800 127.400 145.200 ;
        RECT 127.800 144.800 128.200 145.200 ;
        RECT 129.400 144.800 129.800 145.200 ;
        RECT 125.400 144.100 125.800 144.200 ;
        RECT 126.200 144.100 126.600 144.200 ;
        RECT 125.400 143.800 126.600 144.100 ;
        RECT 128.600 143.800 129.000 144.200 ;
        RECT 118.200 142.800 118.600 143.200 ;
        RECT 124.600 142.800 125.000 143.200 ;
        RECT 127.000 142.800 127.400 143.200 ;
        RECT 116.600 141.800 117.000 142.200 ;
        RECT 118.200 141.800 118.600 142.200 ;
        RECT 123.000 141.800 123.400 142.200 ;
        RECT 126.200 141.800 126.600 142.200 ;
        RECT 115.800 139.800 116.200 140.200 ;
        RECT 111.000 137.800 111.400 138.200 ;
        RECT 113.400 137.800 113.800 138.200 ;
        RECT 111.000 135.200 111.300 137.800 ;
        RECT 113.400 136.200 113.700 137.800 ;
        RECT 113.400 135.800 113.800 136.200 ;
        RECT 111.000 134.800 111.400 135.200 ;
        RECT 114.200 134.800 114.600 135.200 ;
        RECT 110.200 133.800 110.600 134.200 ;
        RECT 110.200 132.200 110.500 133.800 ;
        RECT 107.000 132.100 107.400 132.200 ;
        RECT 107.800 132.100 108.200 132.200 ;
        RECT 107.000 131.800 108.200 132.100 ;
        RECT 110.200 131.800 110.600 132.200 ;
        RECT 108.600 127.800 109.000 128.200 ;
        RECT 109.400 127.800 109.800 128.200 ;
        RECT 110.200 127.800 110.600 128.200 ;
        RECT 108.600 127.200 108.900 127.800 ;
        RECT 109.400 127.200 109.700 127.800 ;
        RECT 110.200 127.200 110.500 127.800 ;
        RECT 107.000 127.100 107.400 127.200 ;
        RECT 107.800 127.100 108.200 127.200 ;
        RECT 107.000 126.800 108.200 127.100 ;
        RECT 108.600 126.800 109.000 127.200 ;
        RECT 109.400 126.800 109.800 127.200 ;
        RECT 110.200 126.800 110.600 127.200 ;
        RECT 111.000 126.200 111.300 134.800 ;
        RECT 112.600 131.800 113.000 132.200 ;
        RECT 112.600 126.200 112.900 131.800 ;
        RECT 107.800 125.800 108.200 126.200 ;
        RECT 110.200 125.800 110.600 126.200 ;
        RECT 111.000 125.800 111.400 126.200 ;
        RECT 111.800 125.800 112.200 126.200 ;
        RECT 112.600 125.800 113.000 126.200 ;
        RECT 113.400 125.800 113.800 126.200 ;
        RECT 107.800 125.200 108.100 125.800 ;
        RECT 106.200 124.800 106.600 125.200 ;
        RECT 107.800 124.800 108.200 125.200 ;
        RECT 106.200 123.200 106.500 124.800 ;
        RECT 106.200 122.800 106.600 123.200 ;
        RECT 107.800 119.200 108.100 124.800 ;
        RECT 110.200 123.200 110.500 125.800 ;
        RECT 110.200 122.800 110.600 123.200 ;
        RECT 111.800 122.200 112.100 125.800 ;
        RECT 113.400 124.200 113.700 125.800 ;
        RECT 113.400 123.800 113.800 124.200 ;
        RECT 111.800 121.800 112.200 122.200 ;
        RECT 114.200 119.200 114.500 134.800 ;
        RECT 115.000 133.800 115.400 134.200 ;
        RECT 115.000 130.200 115.300 133.800 ;
        RECT 115.800 131.800 116.200 132.200 ;
        RECT 115.800 131.200 116.100 131.800 ;
        RECT 115.800 130.800 116.200 131.200 ;
        RECT 115.000 129.800 115.400 130.200 ;
        RECT 115.000 128.200 115.300 129.800 ;
        RECT 115.800 128.800 116.200 129.200 ;
        RECT 115.800 128.200 116.100 128.800 ;
        RECT 115.000 127.800 115.400 128.200 ;
        RECT 115.800 127.800 116.200 128.200 ;
        RECT 116.600 124.200 116.900 141.800 ;
        RECT 118.200 141.200 118.500 141.800 ;
        RECT 123.000 141.200 123.300 141.800 ;
        RECT 118.200 140.800 118.600 141.200 ;
        RECT 123.000 140.800 123.400 141.200 ;
        RECT 118.200 132.100 118.600 137.900 ;
        RECT 119.000 136.800 119.400 137.200 ;
        RECT 119.000 135.200 119.300 136.800 ;
        RECT 119.000 134.800 119.400 135.200 ;
        RECT 121.400 135.000 121.800 135.100 ;
        RECT 122.200 135.000 122.600 135.100 ;
        RECT 121.400 134.700 122.600 135.000 ;
        RECT 123.000 132.100 123.400 137.900 ;
        RECT 126.200 137.200 126.500 141.800 ;
        RECT 125.400 136.800 125.800 137.200 ;
        RECT 126.200 136.800 126.600 137.200 ;
        RECT 125.400 136.200 125.700 136.800 ;
        RECT 123.800 133.800 124.200 134.200 ;
        RECT 117.400 130.800 117.800 131.200 ;
        RECT 117.400 126.200 117.700 130.800 ;
        RECT 118.200 129.800 118.600 130.200 ;
        RECT 118.200 129.200 118.500 129.800 ;
        RECT 118.200 128.800 118.600 129.200 ;
        RECT 117.400 125.800 117.800 126.200 ;
        RECT 116.600 123.800 117.000 124.200 ;
        RECT 119.800 123.800 120.200 124.200 ;
        RECT 116.600 123.100 117.000 123.200 ;
        RECT 117.400 123.100 117.800 123.200 ;
        RECT 116.600 122.800 117.800 123.100 ;
        RECT 107.800 118.800 108.200 119.200 ;
        RECT 108.600 118.800 109.000 119.200 ;
        RECT 114.200 118.800 114.600 119.200 ;
        RECT 105.400 115.800 105.800 116.200 ;
        RECT 106.200 115.800 106.600 116.200 ;
        RECT 105.400 114.200 105.700 115.800 ;
        RECT 106.200 114.200 106.500 115.800 ;
        RECT 107.800 114.800 108.200 115.200 ;
        RECT 107.800 114.200 108.100 114.800 ;
        RECT 108.600 114.200 108.900 118.800 ;
        RECT 119.000 116.800 119.400 117.200 ;
        RECT 109.400 115.800 109.800 116.200 ;
        RECT 113.400 115.900 113.800 116.300 ;
        RECT 116.700 115.900 117.100 116.300 ;
        RECT 109.400 115.200 109.700 115.800 ;
        RECT 109.400 114.800 109.800 115.200 ;
        RECT 113.400 114.200 113.700 115.900 ;
        RECT 115.400 114.200 115.800 114.300 ;
        RECT 105.400 114.100 105.800 114.200 ;
        RECT 104.600 113.800 105.800 114.100 ;
        RECT 106.200 113.800 106.600 114.200 ;
        RECT 107.800 113.800 108.200 114.200 ;
        RECT 108.600 113.800 109.000 114.200 ;
        RECT 111.000 114.100 111.400 114.200 ;
        RECT 111.800 114.100 112.200 114.200 ;
        RECT 111.000 113.800 112.200 114.100 ;
        RECT 112.600 113.800 113.000 114.200 ;
        RECT 113.400 113.900 115.800 114.200 ;
        RECT 104.600 107.200 104.900 113.800 ;
        RECT 104.600 106.800 105.000 107.200 ;
        RECT 102.200 105.800 102.600 106.200 ;
        RECT 103.000 105.800 103.400 106.200 ;
        RECT 103.800 105.800 104.200 106.200 ;
        RECT 102.200 101.200 102.500 105.800 ;
        RECT 103.000 105.200 103.300 105.800 ;
        RECT 103.000 104.800 103.400 105.200 ;
        RECT 102.200 100.800 102.600 101.200 ;
        RECT 102.200 95.200 102.500 100.800 ;
        RECT 102.200 94.800 102.600 95.200 ;
        RECT 103.800 88.200 104.100 105.800 ;
        RECT 104.600 104.100 105.000 104.200 ;
        RECT 105.400 104.100 105.800 104.200 ;
        RECT 104.600 103.800 105.800 104.100 ;
        RECT 107.800 103.100 108.200 108.900 ;
        RECT 104.600 93.100 105.000 95.900 ;
        RECT 105.400 94.800 105.800 95.200 ;
        RECT 105.400 89.200 105.700 94.800 ;
        RECT 106.200 92.100 106.600 97.900 ;
        RECT 107.800 96.800 108.200 97.200 ;
        RECT 107.800 95.200 108.100 96.800 ;
        RECT 108.600 95.200 108.900 113.800 ;
        RECT 112.600 112.200 112.900 113.800 ;
        RECT 113.400 113.500 113.700 113.900 ;
        RECT 114.100 113.500 114.500 113.600 ;
        RECT 115.800 113.500 116.200 113.600 ;
        RECT 116.800 113.500 117.100 115.900 ;
        RECT 119.000 116.200 119.300 116.800 ;
        RECT 119.000 115.800 119.400 116.200 ;
        RECT 117.400 114.100 117.800 114.200 ;
        RECT 118.200 114.100 118.600 114.200 ;
        RECT 117.400 113.800 118.600 114.100 ;
        RECT 113.400 113.100 113.800 113.500 ;
        RECT 114.100 113.200 116.200 113.500 ;
        RECT 116.700 113.100 117.100 113.500 ;
        RECT 112.600 111.800 113.000 112.200 ;
        RECT 115.000 111.800 115.400 112.200 ;
        RECT 110.200 106.100 110.600 106.200 ;
        RECT 111.000 106.100 111.400 106.200 ;
        RECT 110.200 105.800 111.400 106.100 ;
        RECT 112.600 103.100 113.000 108.900 ;
        RECT 113.400 107.800 113.800 108.200 ;
        RECT 113.400 107.200 113.700 107.800 ;
        RECT 113.400 106.800 113.800 107.200 ;
        RECT 114.200 105.100 114.600 107.900 ;
        RECT 115.000 106.200 115.300 111.800 ;
        RECT 119.800 110.100 120.100 123.800 ;
        RECT 120.600 123.100 121.000 128.900 ;
        RECT 123.800 127.200 124.100 133.800 ;
        RECT 124.600 133.100 125.000 135.900 ;
        RECT 125.400 135.800 125.800 136.200 ;
        RECT 127.000 134.200 127.300 142.800 ;
        RECT 127.800 141.800 128.200 142.200 ;
        RECT 127.800 138.200 128.100 141.800 ;
        RECT 128.600 139.200 128.900 143.800 ;
        RECT 128.600 138.800 129.000 139.200 ;
        RECT 127.800 137.800 128.200 138.200 ;
        RECT 129.400 136.200 129.700 144.800 ;
        RECT 131.000 141.800 131.400 142.200 ;
        RECT 131.000 141.200 131.300 141.800 ;
        RECT 131.000 140.800 131.400 141.200 ;
        RECT 131.800 136.200 132.100 145.800 ;
        RECT 135.000 144.200 135.300 145.800 ;
        RECT 135.000 143.800 135.400 144.200 ;
        RECT 138.200 142.200 138.500 146.800 ;
        RECT 139.000 145.100 139.300 146.800 ;
        RECT 141.000 146.700 141.400 146.800 ;
        RECT 142.400 145.100 142.700 147.500 ;
        RECT 139.000 144.700 139.400 145.100 ;
        RECT 142.300 144.700 142.700 145.100 ;
        RECT 143.000 145.100 143.300 148.800 ;
        RECT 146.200 148.200 146.500 151.800 ;
        RECT 152.600 149.200 152.900 153.800 ;
        RECT 153.400 152.100 153.800 157.900 ;
        RECT 154.200 152.100 154.600 158.900 ;
        RECT 155.000 152.100 155.400 158.900 ;
        RECT 158.200 155.800 158.600 156.200 ;
        RECT 158.200 155.200 158.500 155.800 ;
        RECT 158.200 154.800 158.600 155.200 ;
        RECT 159.800 150.200 160.100 166.800 ;
        RECT 160.500 165.100 160.800 167.500 ;
        RECT 161.400 167.400 161.800 167.500 ;
        RECT 163.100 167.400 163.500 167.500 ;
        RECT 163.900 167.100 164.200 167.500 ;
        RECT 161.800 166.800 164.200 167.100 ;
        RECT 161.800 166.700 162.200 166.800 ;
        RECT 161.400 165.800 161.800 166.200 ;
        RECT 160.500 164.700 160.900 165.100 ;
        RECT 161.400 164.200 161.700 165.800 ;
        RECT 163.900 165.100 164.200 166.800 ;
        RECT 163.800 164.700 164.200 165.100 ;
        RECT 164.600 166.800 165.000 167.200 ;
        RECT 164.600 164.200 164.900 166.800 ;
        RECT 165.400 164.200 165.700 171.800 ;
        RECT 167.000 168.800 167.400 169.200 ;
        RECT 167.000 166.200 167.300 168.800 ;
        RECT 167.000 165.800 167.400 166.200 ;
        RECT 161.400 163.800 161.800 164.200 ;
        RECT 164.600 163.800 165.000 164.200 ;
        RECT 165.400 163.800 165.800 164.200 ;
        RECT 169.400 162.100 169.800 168.900 ;
        RECT 170.200 162.100 170.600 168.900 ;
        RECT 171.000 163.100 171.400 168.900 ;
        RECT 171.800 166.800 172.200 167.200 ;
        RECT 171.800 160.200 172.100 166.800 ;
        RECT 172.600 163.100 173.000 168.900 ;
        RECT 173.400 168.200 173.700 172.800 ;
        RECT 173.400 167.800 173.800 168.200 ;
        RECT 171.800 159.800 172.200 160.200 ;
        RECT 162.200 155.100 162.600 155.200 ;
        RECT 163.000 155.100 163.400 155.200 ;
        RECT 162.200 154.800 163.400 155.100 ;
        RECT 165.400 152.100 165.800 158.900 ;
        RECT 166.200 152.100 166.600 158.900 ;
        RECT 167.000 152.100 167.400 157.900 ;
        RECT 167.800 153.800 168.200 154.200 ;
        RECT 167.800 152.200 168.100 153.800 ;
        RECT 167.800 151.800 168.200 152.200 ;
        RECT 168.600 152.100 169.000 157.900 ;
        RECT 169.400 153.800 169.800 154.200 ;
        RECT 169.400 153.200 169.700 153.800 ;
        RECT 169.400 152.800 169.800 153.200 ;
        RECT 170.200 152.100 170.600 157.900 ;
        RECT 171.000 152.100 171.400 158.900 ;
        RECT 171.800 152.100 172.200 158.900 ;
        RECT 172.600 152.100 173.000 158.900 ;
        RECT 173.400 158.200 173.700 167.800 ;
        RECT 174.200 163.100 174.600 168.900 ;
        RECT 175.000 162.100 175.400 168.900 ;
        RECT 175.800 162.100 176.200 168.900 ;
        RECT 176.600 162.100 177.000 168.900 ;
        RECT 177.400 166.200 177.700 174.800 ;
        RECT 178.200 172.100 178.600 178.900 ;
        RECT 179.000 172.100 179.400 178.900 ;
        RECT 179.800 172.100 180.200 177.900 ;
        RECT 180.600 173.800 181.000 174.200 ;
        RECT 180.600 169.200 180.900 173.800 ;
        RECT 181.400 172.100 181.800 177.900 ;
        RECT 182.200 173.800 182.600 174.200 ;
        RECT 182.200 173.200 182.500 173.800 ;
        RECT 182.200 172.800 182.600 173.200 ;
        RECT 183.000 172.100 183.400 177.900 ;
        RECT 183.800 172.100 184.200 178.900 ;
        RECT 184.600 172.100 185.000 178.900 ;
        RECT 185.400 172.100 185.800 178.900 ;
        RECT 195.000 176.800 195.400 177.200 ;
        RECT 195.000 176.200 195.300 176.800 ;
        RECT 195.000 175.800 195.400 176.200 ;
        RECT 194.200 174.800 194.600 175.200 ;
        RECT 192.600 173.100 193.000 173.200 ;
        RECT 193.400 173.100 193.800 173.200 ;
        RECT 192.600 172.800 193.800 173.100 ;
        RECT 190.200 171.800 190.600 172.200 ;
        RECT 191.800 171.800 192.200 172.200 ;
        RECT 190.200 171.200 190.500 171.800 ;
        RECT 190.200 170.800 190.600 171.200 ;
        RECT 180.600 168.800 181.000 169.200 ;
        RECT 184.600 169.100 185.000 169.200 ;
        RECT 185.400 169.100 185.800 169.200 ;
        RECT 184.600 168.800 185.800 169.100 ;
        RECT 190.200 168.800 190.600 169.200 ;
        RECT 190.200 168.200 190.500 168.800 ;
        RECT 187.800 167.800 188.200 168.200 ;
        RECT 190.200 167.800 190.600 168.200 ;
        RECT 191.000 168.100 191.400 168.200 ;
        RECT 191.800 168.100 192.100 171.800 ;
        RECT 194.200 169.200 194.500 174.800 ;
        RECT 195.000 173.800 195.400 174.200 ;
        RECT 195.000 173.200 195.300 173.800 ;
        RECT 195.000 172.800 195.400 173.200 ;
        RECT 196.600 172.800 197.000 173.200 ;
        RECT 200.600 173.100 201.000 173.200 ;
        RECT 201.400 173.100 201.800 173.200 ;
        RECT 200.600 172.800 201.800 173.100 ;
        RECT 202.200 172.800 202.600 173.200 ;
        RECT 196.600 172.200 196.900 172.800 ;
        RECT 196.600 171.800 197.000 172.200 ;
        RECT 194.200 168.800 194.600 169.200 ;
        RECT 191.000 167.800 192.100 168.100 ;
        RECT 192.700 167.800 193.100 167.900 ;
        RECT 187.800 167.200 188.100 167.800 ;
        RECT 192.700 167.500 195.500 167.800 ;
        RECT 195.800 167.500 196.200 167.900 ;
        RECT 183.000 167.100 183.400 167.200 ;
        RECT 183.800 167.100 184.200 167.200 ;
        RECT 183.000 166.800 184.200 167.100 ;
        RECT 187.800 166.800 188.200 167.200 ;
        RECT 189.400 166.800 189.800 167.200 ;
        RECT 191.000 167.100 191.400 167.200 ;
        RECT 191.800 167.100 192.200 167.200 ;
        RECT 191.000 166.800 192.200 167.100 ;
        RECT 189.400 166.200 189.700 166.800 ;
        RECT 177.400 165.800 177.800 166.200 ;
        RECT 187.000 165.800 187.400 166.200 ;
        RECT 188.600 165.800 189.000 166.200 ;
        RECT 189.400 165.800 189.800 166.200 ;
        RECT 187.000 165.200 187.300 165.800 ;
        RECT 179.800 164.800 180.200 165.200 ;
        RECT 183.800 165.100 184.200 165.200 ;
        RECT 184.600 165.100 185.000 165.200 ;
        RECT 183.800 164.800 185.000 165.100 ;
        RECT 187.000 164.800 187.400 165.200 ;
        RECT 179.800 159.200 180.100 164.800 ;
        RECT 181.400 161.800 181.800 162.200 ;
        RECT 179.800 158.800 180.200 159.200 ;
        RECT 173.400 157.800 173.800 158.200 ;
        RECT 173.400 153.200 173.700 157.800 ;
        RECT 179.000 155.800 179.400 156.200 ;
        RECT 179.000 155.200 179.300 155.800 ;
        RECT 179.000 155.100 179.400 155.200 ;
        RECT 178.200 154.800 179.400 155.100 ;
        RECT 180.600 154.800 181.000 155.200 ;
        RECT 173.400 152.800 173.800 153.200 ;
        RECT 177.400 152.100 177.800 152.200 ;
        RECT 176.600 151.800 177.800 152.100 ;
        RECT 159.800 149.800 160.200 150.200 ;
        RECT 163.000 149.800 163.400 150.200 ;
        RECT 152.600 148.800 153.000 149.200 ;
        RECT 154.200 149.100 154.600 149.200 ;
        RECT 155.000 149.100 155.400 149.200 ;
        RECT 154.200 148.800 155.400 149.100 ;
        RECT 146.200 147.800 146.600 148.200 ;
        RECT 151.000 148.100 151.400 148.200 ;
        RECT 151.800 148.100 152.200 148.200 ;
        RECT 151.000 147.800 152.200 148.100 ;
        RECT 146.200 147.200 146.500 147.800 ;
        RECT 159.800 147.200 160.100 149.800 ;
        RECT 160.600 148.100 161.000 148.200 ;
        RECT 161.400 148.100 161.800 148.200 ;
        RECT 160.600 147.800 161.800 148.100 ;
        RECT 143.800 146.800 144.200 147.200 ;
        RECT 146.200 146.800 146.600 147.200 ;
        RECT 149.400 146.800 149.800 147.200 ;
        RECT 154.200 147.100 154.600 147.200 ;
        RECT 154.200 146.800 155.300 147.100 ;
        RECT 143.800 146.200 144.100 146.800 ;
        RECT 143.800 145.800 144.200 146.200 ;
        RECT 148.600 145.800 149.000 146.200 ;
        RECT 143.000 144.800 144.100 145.100 ;
        RECT 142.200 143.800 142.600 144.200 ;
        RECT 138.200 141.800 138.600 142.200 ;
        RECT 141.400 139.800 141.800 140.200 ;
        RECT 141.400 139.200 141.700 139.800 ;
        RECT 141.400 138.800 141.800 139.200 ;
        RECT 140.600 137.800 141.000 138.200 ;
        RECT 129.400 135.800 129.800 136.200 ;
        RECT 131.800 135.800 132.200 136.200 ;
        RECT 134.200 135.800 134.600 136.200 ;
        RECT 131.800 135.200 132.100 135.800 ;
        RECT 134.200 135.200 134.500 135.800 ;
        RECT 130.200 135.100 130.600 135.200 ;
        RECT 131.000 135.100 131.400 135.200 ;
        RECT 130.200 134.800 131.400 135.100 ;
        RECT 131.800 134.800 132.200 135.200 ;
        RECT 134.200 134.800 134.600 135.200 ;
        RECT 135.800 135.100 136.200 135.200 ;
        RECT 136.600 135.100 137.000 135.200 ;
        RECT 135.800 134.800 137.000 135.100 ;
        RECT 137.400 135.100 137.800 135.200 ;
        RECT 138.200 135.100 138.600 135.200 ;
        RECT 137.400 134.800 138.600 135.100 ;
        RECT 139.800 134.800 140.200 135.200 ;
        RECT 127.000 133.800 127.400 134.200 ;
        RECT 134.200 133.800 134.600 134.200 ;
        RECT 134.200 133.200 134.500 133.800 ;
        RECT 125.400 133.100 125.800 133.200 ;
        RECT 126.200 133.100 126.600 133.200 ;
        RECT 125.400 132.800 126.600 133.100 ;
        RECT 131.800 133.100 132.200 133.200 ;
        RECT 132.600 133.100 133.000 133.200 ;
        RECT 131.800 132.800 133.000 133.100 ;
        RECT 134.200 132.800 134.600 133.200 ;
        RECT 135.000 132.800 135.400 133.200 ;
        RECT 135.000 131.200 135.300 132.800 ;
        RECT 135.000 130.800 135.400 131.200 ;
        RECT 123.800 126.800 124.200 127.200 ;
        RECT 123.000 126.100 123.400 126.200 ;
        RECT 123.800 126.100 124.200 126.200 ;
        RECT 123.000 125.800 124.200 126.100 ;
        RECT 122.200 123.800 122.600 124.200 ;
        RECT 120.600 116.100 121.000 116.200 ;
        RECT 121.400 116.100 121.800 116.200 ;
        RECT 120.600 115.800 121.800 116.100 ;
        RECT 120.600 114.800 121.000 115.200 ;
        RECT 120.600 112.200 120.900 114.800 ;
        RECT 120.600 111.800 121.000 112.200 ;
        RECT 119.800 109.800 120.900 110.100 ;
        RECT 115.000 105.800 115.400 106.200 ;
        RECT 114.200 102.800 114.600 103.200 ;
        RECT 107.800 94.800 108.200 95.200 ;
        RECT 108.600 94.800 109.000 95.200 ;
        RECT 110.200 94.800 110.600 95.200 ;
        RECT 105.400 88.800 105.800 89.200 ;
        RECT 100.600 87.800 101.000 88.200 ;
        RECT 103.800 87.800 104.200 88.200 ;
        RECT 105.400 87.200 105.700 88.800 ;
        RECT 103.000 86.800 103.400 87.200 ;
        RECT 105.400 86.800 105.800 87.200 ;
        RECT 106.200 86.800 106.600 87.200 ;
        RECT 100.600 85.800 101.000 86.200 ;
        RECT 100.600 85.200 100.900 85.800 ;
        RECT 103.000 85.200 103.300 86.800 ;
        RECT 106.200 86.200 106.500 86.800 ;
        RECT 103.800 86.100 104.200 86.200 ;
        RECT 104.600 86.100 105.000 86.200 ;
        RECT 103.800 85.800 105.000 86.100 ;
        RECT 106.200 85.800 106.600 86.200 ;
        RECT 100.600 84.800 101.000 85.200 ;
        RECT 103.000 84.800 103.400 85.200 ;
        RECT 95.800 76.800 96.200 77.200 ;
        RECT 97.400 75.800 97.800 76.200 ;
        RECT 95.800 75.100 96.200 75.200 ;
        RECT 96.600 75.100 97.000 75.200 ;
        RECT 95.800 74.800 97.000 75.100 ;
        RECT 97.400 74.200 97.700 75.800 ;
        RECT 97.400 74.100 97.800 74.200 ;
        RECT 98.200 74.100 98.600 74.200 ;
        RECT 97.400 73.800 98.600 74.100 ;
        RECT 94.200 72.800 94.600 73.200 ;
        RECT 95.000 73.100 95.400 73.200 ;
        RECT 95.800 73.100 96.200 73.200 ;
        RECT 95.000 72.800 96.200 73.100 ;
        RECT 99.000 72.100 99.400 77.900 ;
        RECT 99.800 77.800 100.200 78.200 ;
        RECT 102.200 74.800 102.600 75.200 ;
        RECT 99.800 73.800 100.200 74.200 ;
        RECT 93.400 68.800 93.800 69.200 ;
        RECT 99.000 68.800 99.400 69.200 ;
        RECT 99.000 68.200 99.300 68.800 ;
        RECT 99.000 67.800 99.400 68.200 ;
        RECT 92.600 67.100 93.000 67.200 ;
        RECT 93.400 67.100 93.800 67.200 ;
        RECT 92.600 66.800 93.800 67.100 ;
        RECT 98.200 67.100 98.600 67.200 ;
        RECT 99.000 67.100 99.400 67.200 ;
        RECT 98.200 66.800 99.400 67.100 ;
        RECT 84.600 65.800 85.700 66.100 ;
        RECT 86.200 65.800 86.600 66.200 ;
        RECT 90.200 65.800 90.600 66.200 ;
        RECT 91.800 65.800 92.200 66.200 ;
        RECT 93.400 65.800 93.800 66.200 ;
        RECT 83.800 64.800 84.200 65.200 ;
        RECT 84.600 64.800 85.000 65.200 ;
        RECT 83.000 56.800 83.400 57.200 ;
        RECT 83.800 54.200 84.100 64.800 ;
        RECT 84.600 64.200 84.900 64.800 ;
        RECT 86.200 64.200 86.500 65.800 ;
        RECT 90.200 65.200 90.500 65.800 ;
        RECT 93.400 65.200 93.700 65.800 ;
        RECT 87.800 64.800 88.200 65.200 ;
        RECT 90.200 64.800 90.600 65.200 ;
        RECT 93.400 64.800 93.800 65.200 ;
        RECT 95.800 65.100 96.200 65.200 ;
        RECT 96.600 65.100 97.000 65.200 ;
        RECT 95.800 64.800 97.000 65.100 ;
        RECT 84.600 64.100 85.000 64.200 ;
        RECT 84.600 63.800 85.700 64.100 ;
        RECT 86.200 63.800 86.600 64.200 ;
        RECT 85.400 63.200 85.700 63.800 ;
        RECT 85.400 62.800 85.800 63.200 ;
        RECT 84.600 56.800 85.000 57.200 ;
        RECT 84.600 55.200 84.900 56.800 ;
        RECT 85.400 56.200 85.700 62.800 ;
        RECT 87.800 62.200 88.100 64.800 ;
        RECT 87.800 61.800 88.200 62.200 ;
        RECT 88.600 60.800 89.000 61.200 ;
        RECT 87.000 59.800 87.400 60.200 ;
        RECT 87.000 59.200 87.300 59.800 ;
        RECT 87.000 58.800 87.400 59.200 ;
        RECT 85.400 55.800 85.800 56.200 ;
        RECT 84.600 54.800 85.000 55.200 ;
        RECT 87.000 54.800 87.400 55.200 ;
        RECT 81.400 53.800 81.800 54.200 ;
        RECT 83.800 53.800 84.200 54.200 ;
        RECT 77.400 46.800 77.800 47.200 ;
        RECT 75.000 40.800 75.400 41.200 ;
        RECT 73.400 39.800 73.800 40.200 ;
        RECT 73.400 35.200 73.700 39.800 ;
        RECT 75.000 39.200 75.300 40.800 ;
        RECT 79.800 39.200 80.100 53.800 ;
        RECT 82.200 53.100 82.600 53.200 ;
        RECT 81.400 52.800 82.600 53.100 ;
        RECT 83.000 52.800 83.400 53.200 ;
        RECT 80.600 46.800 81.000 47.200 ;
        RECT 80.600 46.200 80.900 46.800 ;
        RECT 80.600 45.800 81.000 46.200 ;
        RECT 75.000 38.800 75.400 39.200 ;
        RECT 79.800 38.800 80.200 39.200 ;
        RECT 80.600 36.800 81.000 37.200 ;
        RECT 80.600 36.200 80.900 36.800 ;
        RECT 75.000 35.800 75.400 36.200 ;
        RECT 80.600 35.800 81.000 36.200 ;
        RECT 73.400 34.800 73.800 35.200 ;
        RECT 70.200 34.100 70.600 34.200 ;
        RECT 69.400 33.800 70.600 34.100 ;
        RECT 53.400 33.200 53.700 33.800 ;
        RECT 58.200 33.200 58.500 33.800 ;
        RECT 53.400 32.800 53.800 33.200 ;
        RECT 54.200 32.800 54.600 33.200 ;
        RECT 56.600 32.800 57.000 33.200 ;
        RECT 57.400 32.800 57.800 33.200 ;
        RECT 58.200 32.800 58.600 33.200 ;
        RECT 54.200 31.200 54.500 32.800 ;
        RECT 54.200 30.800 54.600 31.200 ;
        RECT 55.000 29.800 55.400 30.200 ;
        RECT 55.000 27.200 55.300 29.800 ;
        RECT 55.000 26.800 55.400 27.200 ;
        RECT 55.800 26.800 56.200 27.200 ;
        RECT 55.800 26.200 56.100 26.800 ;
        RECT 54.200 26.100 54.600 26.200 ;
        RECT 55.000 26.100 55.400 26.200 ;
        RECT 54.200 25.800 55.400 26.100 ;
        RECT 55.800 25.800 56.200 26.200 ;
        RECT 56.600 18.200 56.900 32.800 ;
        RECT 57.400 25.200 57.700 32.800 ;
        RECT 59.000 30.800 59.400 31.200 ;
        RECT 59.000 29.200 59.300 30.800 ;
        RECT 61.400 30.200 61.700 33.800 ;
        RECT 61.400 30.100 61.800 30.200 ;
        RECT 60.600 29.800 61.800 30.100 ;
        RECT 59.000 28.800 59.400 29.200 ;
        RECT 59.800 26.800 60.200 27.200 ;
        RECT 59.000 25.800 59.400 26.200 ;
        RECT 57.400 24.800 57.800 25.200 ;
        RECT 59.000 19.200 59.300 25.800 ;
        RECT 59.800 23.200 60.100 26.800 ;
        RECT 60.600 26.200 60.900 29.800 ;
        RECT 61.400 27.800 61.800 28.200 ;
        RECT 61.400 27.200 61.700 27.800 ;
        RECT 61.400 26.800 61.800 27.200 ;
        RECT 60.600 25.800 61.000 26.200 ;
        RECT 62.200 26.100 62.500 33.800 ;
        RECT 69.400 31.800 69.800 32.200 ;
        RECT 71.800 31.800 72.200 32.200 ;
        RECT 67.000 29.800 67.400 30.200 ;
        RECT 63.000 27.800 63.400 28.200 ;
        RECT 63.000 27.200 63.300 27.800 ;
        RECT 67.000 27.200 67.300 29.800 ;
        RECT 69.400 29.200 69.700 31.800 ;
        RECT 71.800 30.200 72.100 31.800 ;
        RECT 71.800 29.800 72.200 30.200 ;
        RECT 75.000 29.200 75.300 35.800 ;
        RECT 81.400 35.200 81.700 52.800 ;
        RECT 83.000 52.200 83.300 52.800 ;
        RECT 83.000 51.800 83.400 52.200 ;
        RECT 83.800 51.800 84.200 52.200 ;
        RECT 83.800 51.200 84.100 51.800 ;
        RECT 84.600 51.200 84.900 54.800 ;
        RECT 87.000 53.200 87.300 54.800 ;
        RECT 88.600 54.200 88.900 60.800 ;
        RECT 98.200 59.800 98.600 60.200 ;
        RECT 89.400 55.800 89.800 56.200 ;
        RECT 91.000 56.100 91.400 56.200 ;
        RECT 91.800 56.100 92.200 56.200 ;
        RECT 91.000 55.800 92.200 56.100 ;
        RECT 92.600 55.800 93.000 56.200 ;
        RECT 89.400 55.200 89.700 55.800 ;
        RECT 89.400 54.800 89.800 55.200 ;
        RECT 92.600 55.100 92.900 55.800 ;
        RECT 91.800 54.800 92.900 55.100 ;
        RECT 91.800 54.200 92.100 54.800 ;
        RECT 87.800 53.800 88.200 54.200 ;
        RECT 88.600 53.800 89.000 54.200 ;
        RECT 91.800 53.800 92.200 54.200 ;
        RECT 93.400 53.800 93.800 54.200 ;
        RECT 87.800 53.200 88.100 53.800 ;
        RECT 93.400 53.200 93.700 53.800 ;
        RECT 87.000 52.800 87.400 53.200 ;
        RECT 87.800 52.800 88.200 53.200 ;
        RECT 90.200 52.800 90.600 53.200 ;
        RECT 93.400 52.800 93.800 53.200 ;
        RECT 94.200 53.100 94.600 55.900 ;
        RECT 83.800 50.800 84.200 51.200 ;
        RECT 84.600 50.800 85.000 51.200 ;
        RECT 88.600 50.800 89.000 51.200 ;
        RECT 82.200 47.800 82.600 48.200 ;
        RECT 83.000 47.800 83.400 48.200 ;
        RECT 82.200 47.200 82.500 47.800 ;
        RECT 82.200 46.800 82.600 47.200 ;
        RECT 82.200 45.800 82.600 46.200 ;
        RECT 82.200 45.200 82.500 45.800 ;
        RECT 82.200 44.800 82.600 45.200 ;
        RECT 82.200 41.200 82.500 44.800 ;
        RECT 82.200 40.800 82.600 41.200 ;
        RECT 83.000 40.200 83.300 47.800 ;
        RECT 83.000 39.800 83.400 40.200 ;
        RECT 77.400 34.800 77.800 35.200 ;
        RECT 79.800 34.800 80.200 35.200 ;
        RECT 81.400 34.800 81.800 35.200 ;
        RECT 82.200 34.800 82.600 35.200 ;
        RECT 77.400 34.200 77.700 34.800 ;
        RECT 77.400 33.800 77.800 34.200 ;
        RECT 79.800 33.200 80.100 34.800 ;
        RECT 75.800 32.800 76.200 33.200 ;
        RECT 78.200 32.800 78.600 33.200 ;
        RECT 79.800 32.800 80.200 33.200 ;
        RECT 69.400 28.800 69.800 29.200 ;
        RECT 75.000 28.800 75.400 29.200 ;
        RECT 63.000 26.800 63.400 27.200 ;
        RECT 65.400 27.100 65.800 27.200 ;
        RECT 66.200 27.100 66.600 27.200 ;
        RECT 65.400 26.800 66.600 27.100 ;
        RECT 67.000 26.800 67.400 27.200 ;
        RECT 69.400 26.800 69.800 27.200 ;
        RECT 71.800 27.100 72.200 27.200 ;
        RECT 72.600 27.100 73.000 27.200 ;
        RECT 71.800 26.800 73.000 27.100 ;
        RECT 63.000 26.100 63.400 26.200 ;
        RECT 62.200 25.800 63.400 26.100 ;
        RECT 66.200 25.800 66.600 26.200 ;
        RECT 67.800 25.800 68.200 26.200 ;
        RECT 62.200 23.200 62.500 25.800 ;
        RECT 63.000 25.100 63.400 25.200 ;
        RECT 63.800 25.100 64.200 25.200 ;
        RECT 63.000 24.800 64.200 25.100 ;
        RECT 65.400 24.800 65.800 25.200 ;
        RECT 65.400 24.200 65.700 24.800 ;
        RECT 65.400 23.800 65.800 24.200 ;
        RECT 59.800 22.800 60.200 23.200 ;
        RECT 60.600 22.800 61.000 23.200 ;
        RECT 62.200 22.800 62.600 23.200 ;
        RECT 59.000 18.800 59.400 19.200 ;
        RECT 56.600 17.800 57.000 18.200 ;
        RECT 55.000 16.800 55.400 17.200 ;
        RECT 55.000 16.200 55.300 16.800 ;
        RECT 55.000 15.800 55.400 16.200 ;
        RECT 52.600 14.800 53.000 15.200 ;
        RECT 53.400 14.800 53.800 15.200 ;
        RECT 53.400 14.200 53.700 14.800 ;
        RECT 56.600 14.200 56.900 17.800 ;
        RECT 59.800 15.100 60.200 15.200 ;
        RECT 60.600 15.100 60.900 22.800 ;
        RECT 66.200 22.200 66.500 25.800 ;
        RECT 62.200 21.800 62.600 22.200 ;
        RECT 66.200 21.800 66.600 22.200 ;
        RECT 62.200 19.200 62.500 21.800 ;
        RECT 67.800 19.200 68.100 25.800 ;
        RECT 69.400 25.200 69.700 26.800 ;
        RECT 72.600 26.100 73.000 26.200 ;
        RECT 73.400 26.100 73.800 26.200 ;
        RECT 72.600 25.800 73.800 26.100 ;
        RECT 74.200 25.800 74.600 26.200 ;
        RECT 74.200 25.200 74.500 25.800 ;
        RECT 69.400 24.800 69.800 25.200 ;
        RECT 70.200 24.800 70.600 25.200 ;
        RECT 71.800 25.100 72.200 25.200 ;
        RECT 72.600 25.100 73.000 25.200 ;
        RECT 71.800 24.800 73.000 25.100 ;
        RECT 74.200 24.800 74.600 25.200 ;
        RECT 68.600 22.800 69.000 23.200 ;
        RECT 62.200 18.800 62.600 19.200 ;
        RECT 67.800 18.800 68.200 19.200 ;
        RECT 59.800 14.800 60.900 15.100 ;
        RECT 61.400 14.800 61.800 15.200 ;
        RECT 61.400 14.200 61.700 14.800 ;
        RECT 51.800 13.800 52.200 14.200 ;
        RECT 53.400 13.800 53.800 14.200 ;
        RECT 56.600 13.800 57.000 14.200 ;
        RECT 61.400 13.800 61.800 14.200 ;
        RECT 57.400 12.800 57.800 13.200 ;
        RECT 61.400 12.800 61.800 13.200 ;
        RECT 57.400 12.200 57.700 12.800 ;
        RECT 57.400 11.800 57.800 12.200 ;
        RECT 41.400 5.800 41.800 6.200 ;
        RECT 43.800 5.800 44.200 6.200 ;
        RECT 39.800 4.800 40.200 5.200 ;
        RECT 41.400 4.800 41.800 5.200 ;
        RECT 41.400 4.200 41.700 4.800 ;
        RECT 41.400 3.800 41.800 4.200 ;
        RECT 45.400 3.100 45.800 8.900 ;
        RECT 46.200 6.100 46.600 6.200 ;
        RECT 47.000 6.100 47.400 6.200 ;
        RECT 46.200 5.800 47.400 6.100 ;
        RECT 48.600 5.800 49.000 6.200 ;
        RECT 48.600 5.200 48.900 5.800 ;
        RECT 48.600 4.800 49.000 5.200 ;
        RECT 50.200 3.100 50.600 8.900 ;
        RECT 51.800 5.100 52.200 7.900 ;
        RECT 54.200 5.100 54.600 7.900 ;
        RECT 55.800 3.100 56.200 8.900 ;
        RECT 59.800 7.800 60.200 8.200 ;
        RECT 59.800 7.200 60.100 7.800 ;
        RECT 59.800 6.800 60.200 7.200 ;
        RECT 57.400 6.100 57.800 6.200 ;
        RECT 58.200 6.100 58.600 6.200 ;
        RECT 57.400 5.800 58.600 6.100 ;
        RECT 60.600 3.100 61.000 8.900 ;
        RECT 61.400 8.200 61.700 12.800 ;
        RECT 64.600 12.100 65.000 17.900 ;
        RECT 67.800 16.800 68.200 17.200 ;
        RECT 61.400 7.800 61.800 8.200 ;
        RECT 65.400 6.800 65.800 7.200 ;
        RECT 65.400 6.200 65.700 6.800 ;
        RECT 67.800 6.200 68.100 16.800 ;
        RECT 68.600 15.100 68.900 22.800 ;
        RECT 69.400 19.200 69.700 24.800 ;
        RECT 70.200 24.200 70.500 24.800 ;
        RECT 70.200 23.800 70.600 24.200 ;
        RECT 69.400 18.800 69.800 19.200 ;
        RECT 68.600 14.700 69.000 15.100 ;
        RECT 69.400 12.100 69.800 17.900 ;
        RECT 72.600 16.800 73.000 17.200 ;
        RECT 70.200 13.800 70.600 14.200 ;
        RECT 68.600 10.800 69.000 11.200 ;
        RECT 68.600 8.200 68.900 10.800 ;
        RECT 70.200 8.200 70.500 13.800 ;
        RECT 71.000 13.100 71.400 15.900 ;
        RECT 72.600 15.200 72.900 16.800 ;
        RECT 74.200 15.800 74.600 16.200 ;
        RECT 75.800 16.100 76.100 32.800 ;
        RECT 78.200 32.200 78.500 32.800 ;
        RECT 82.200 32.200 82.500 34.800 ;
        RECT 83.800 34.200 84.100 50.800 ;
        RECT 87.000 49.800 87.400 50.200 ;
        RECT 87.000 49.200 87.300 49.800 ;
        RECT 87.000 48.800 87.400 49.200 ;
        RECT 87.800 48.800 88.200 49.200 ;
        RECT 87.800 48.200 88.100 48.800 ;
        RECT 87.800 47.800 88.200 48.200 ;
        RECT 84.600 46.800 85.000 47.200 ;
        RECT 84.600 46.200 84.900 46.800 ;
        RECT 88.600 46.200 88.900 50.800 ;
        RECT 90.200 49.200 90.500 52.800 ;
        RECT 95.800 52.100 96.200 57.900 ;
        RECT 96.600 55.800 97.000 56.200 ;
        RECT 96.600 55.100 96.900 55.800 ;
        RECT 96.600 54.700 97.000 55.100 ;
        RECT 91.800 50.800 92.200 51.200 ;
        RECT 90.200 48.800 90.600 49.200 ;
        RECT 91.000 48.800 91.400 49.200 ;
        RECT 91.000 48.200 91.300 48.800 ;
        RECT 91.000 47.800 91.400 48.200 ;
        RECT 91.800 47.200 92.100 50.800 ;
        RECT 95.800 49.800 96.200 50.200 ;
        RECT 94.200 49.100 94.600 49.200 ;
        RECT 95.000 49.100 95.400 49.200 ;
        RECT 94.200 48.800 95.400 49.100 ;
        RECT 95.800 47.200 96.100 49.800 ;
        RECT 89.400 46.800 89.800 47.200 ;
        RECT 91.800 46.800 92.200 47.200 ;
        RECT 92.600 46.800 93.000 47.200 ;
        RECT 95.000 46.800 95.400 47.200 ;
        RECT 95.800 46.800 96.200 47.200 ;
        RECT 97.400 46.800 97.800 47.200 ;
        RECT 84.600 45.800 85.000 46.200 ;
        RECT 85.400 45.800 85.800 46.200 ;
        RECT 86.200 45.800 86.600 46.200 ;
        RECT 88.600 45.800 89.000 46.200 ;
        RECT 84.600 38.800 85.000 39.200 ;
        RECT 84.600 35.200 84.900 38.800 ;
        RECT 85.400 37.200 85.700 45.800 ;
        RECT 86.200 45.200 86.500 45.800 ;
        RECT 86.200 44.800 86.600 45.200 ;
        RECT 89.400 43.200 89.700 46.800 ;
        RECT 92.600 46.200 92.900 46.800 ;
        RECT 92.600 45.800 93.000 46.200 ;
        RECT 95.000 45.200 95.300 46.800 ;
        RECT 97.400 46.200 97.700 46.800 ;
        RECT 98.200 46.200 98.500 59.800 ;
        RECT 99.800 55.200 100.100 73.800 ;
        RECT 102.200 73.200 102.500 74.800 ;
        RECT 102.200 72.800 102.600 73.200 ;
        RECT 103.800 72.100 104.200 77.900 ;
        RECT 104.600 76.200 104.900 85.800 ;
        RECT 108.600 83.100 109.000 88.900 ;
        RECT 110.200 87.200 110.500 94.800 ;
        RECT 111.000 92.100 111.400 97.900 ;
        RECT 113.400 96.800 113.800 97.200 ;
        RECT 113.400 95.200 113.700 96.800 ;
        RECT 113.400 94.800 113.800 95.200 ;
        RECT 114.200 94.200 114.500 102.800 ;
        RECT 115.000 98.200 115.300 105.800 ;
        RECT 118.200 105.100 118.600 107.900 ;
        RECT 116.600 103.100 117.000 103.200 ;
        RECT 117.400 103.100 117.800 103.200 ;
        RECT 119.800 103.100 120.200 108.900 ;
        RECT 120.600 108.200 120.900 109.800 ;
        RECT 121.400 108.800 121.800 109.200 ;
        RECT 120.600 107.800 121.000 108.200 ;
        RECT 120.600 107.200 120.900 107.800 ;
        RECT 120.600 106.800 121.000 107.200 ;
        RECT 121.400 106.200 121.700 108.800 ;
        RECT 121.400 105.800 121.800 106.200 ;
        RECT 116.600 102.800 117.800 103.100 ;
        RECT 115.000 97.800 115.400 98.200 ;
        RECT 116.600 97.800 117.000 98.200 ;
        RECT 116.600 96.200 116.900 97.800 ;
        RECT 118.200 96.800 118.600 97.200 ;
        RECT 116.600 95.800 117.000 96.200 ;
        RECT 115.000 95.100 115.400 95.200 ;
        RECT 115.800 95.100 116.200 95.200 ;
        RECT 115.000 94.800 116.200 95.100 ;
        RECT 112.600 93.800 113.000 94.200 ;
        RECT 114.200 93.800 114.600 94.200 ;
        RECT 115.800 93.800 116.200 94.200 ;
        RECT 110.200 86.800 110.600 87.200 ;
        RECT 110.200 85.800 110.600 86.200 ;
        RECT 110.200 85.200 110.500 85.800 ;
        RECT 110.200 84.800 110.600 85.200 ;
        RECT 104.600 75.800 105.000 76.200 ;
        RECT 108.600 76.100 109.000 76.200 ;
        RECT 109.400 76.100 109.800 76.200 ;
        RECT 104.600 73.800 105.000 74.200 ;
        RECT 103.000 66.800 103.400 67.200 ;
        RECT 101.400 65.800 101.800 66.200 ;
        RECT 102.200 65.800 102.600 66.200 ;
        RECT 101.400 58.200 101.700 65.800 ;
        RECT 102.200 65.200 102.500 65.800 ;
        RECT 102.200 64.800 102.600 65.200 ;
        RECT 99.800 54.800 100.200 55.200 ;
        RECT 95.800 46.100 96.200 46.200 ;
        RECT 96.600 46.100 97.000 46.200 ;
        RECT 95.800 45.800 97.000 46.100 ;
        RECT 97.400 45.800 97.800 46.200 ;
        RECT 98.200 45.800 98.600 46.200 ;
        RECT 93.400 45.100 93.800 45.200 ;
        RECT 94.200 45.100 94.600 45.200 ;
        RECT 93.400 44.800 94.600 45.100 ;
        RECT 95.000 44.800 95.400 45.200 ;
        RECT 98.200 44.200 98.500 45.800 ;
        RECT 98.200 43.800 98.600 44.200 ;
        RECT 89.400 42.800 89.800 43.200 ;
        RECT 89.400 39.800 89.800 40.200 ;
        RECT 89.400 39.200 89.700 39.800 ;
        RECT 87.000 38.800 87.400 39.200 ;
        RECT 89.400 38.800 89.800 39.200 ;
        RECT 85.400 36.800 85.800 37.200 ;
        RECT 84.600 34.800 85.000 35.200 ;
        RECT 83.000 33.800 83.400 34.200 ;
        RECT 83.800 33.800 84.200 34.200 ;
        RECT 78.200 31.800 78.600 32.200 ;
        RECT 80.600 31.800 81.000 32.200 ;
        RECT 82.200 31.800 82.600 32.200 ;
        RECT 77.400 29.800 77.800 30.200 ;
        RECT 76.600 26.800 77.000 27.200 ;
        RECT 76.600 26.200 76.900 26.800 ;
        RECT 77.400 26.200 77.700 29.800 ;
        RECT 78.200 26.800 78.600 27.200 ;
        RECT 79.800 26.800 80.200 27.200 ;
        RECT 76.600 25.800 77.000 26.200 ;
        RECT 77.400 25.800 77.800 26.200 ;
        RECT 75.000 15.800 76.100 16.100 ;
        RECT 77.400 23.800 77.800 24.200 ;
        RECT 77.400 16.200 77.700 23.800 ;
        RECT 78.200 22.200 78.500 26.800 ;
        RECT 79.800 25.200 80.100 26.800 ;
        RECT 79.800 24.800 80.200 25.200 ;
        RECT 78.200 21.800 78.600 22.200 ;
        RECT 79.800 20.800 80.200 21.200 ;
        RECT 79.800 19.200 80.100 20.800 ;
        RECT 79.800 18.800 80.200 19.200 ;
        RECT 77.400 15.800 77.800 16.200 ;
        RECT 72.600 14.800 73.000 15.200 ;
        RECT 71.800 14.100 72.200 14.200 ;
        RECT 72.600 14.100 73.000 14.200 ;
        RECT 71.800 13.800 73.000 14.100 ;
        RECT 74.200 13.200 74.500 15.800 ;
        RECT 75.000 14.200 75.300 15.800 ;
        RECT 75.800 14.800 76.200 15.200 ;
        RECT 79.000 15.100 79.400 15.200 ;
        RECT 79.800 15.100 80.200 15.200 ;
        RECT 79.000 14.800 80.200 15.100 ;
        RECT 75.000 13.800 75.400 14.200 ;
        RECT 74.200 12.800 74.600 13.200 ;
        RECT 74.200 11.800 74.600 12.200 ;
        RECT 68.600 7.800 69.000 8.200 ;
        RECT 68.600 7.200 68.900 7.800 ;
        RECT 68.600 6.800 69.000 7.200 ;
        RECT 65.400 5.800 65.800 6.200 ;
        RECT 67.800 5.800 68.200 6.200 ;
        RECT 67.800 5.200 68.100 5.800 ;
        RECT 65.400 5.100 65.800 5.200 ;
        RECT 66.200 5.100 66.600 5.200 ;
        RECT 65.400 4.800 66.600 5.100 ;
        RECT 67.800 4.800 68.200 5.200 ;
        RECT 69.400 5.100 69.800 7.900 ;
        RECT 70.200 7.800 70.600 8.200 ;
        RECT 70.200 7.200 70.500 7.800 ;
        RECT 70.200 6.800 70.600 7.200 ;
        RECT 71.000 3.100 71.400 8.900 ;
        RECT 74.200 6.200 74.500 11.800 ;
        RECT 75.800 10.200 76.100 14.800 ;
        RECT 79.000 12.800 79.400 13.200 ;
        RECT 75.800 9.800 76.200 10.200 ;
        RECT 79.000 9.200 79.300 12.800 ;
        RECT 74.200 5.800 74.600 6.200 ;
        RECT 75.800 3.100 76.200 8.900 ;
        RECT 78.200 8.800 78.600 9.200 ;
        RECT 79.000 8.800 79.400 9.200 ;
        RECT 78.200 8.200 78.500 8.800 ;
        RECT 80.600 8.200 80.900 31.800 ;
        RECT 83.000 30.200 83.300 33.800 ;
        RECT 83.000 30.100 83.400 30.200 ;
        RECT 83.000 29.800 84.100 30.100 ;
        RECT 82.200 28.800 82.600 29.200 ;
        RECT 82.200 26.200 82.500 28.800 ;
        RECT 83.000 27.800 83.400 28.200 ;
        RECT 83.000 27.200 83.300 27.800 ;
        RECT 83.800 27.200 84.100 29.800 ;
        RECT 84.600 27.200 84.900 34.800 ;
        RECT 85.400 28.200 85.700 36.800 ;
        RECT 87.000 36.200 87.300 38.800 ;
        RECT 87.000 35.800 87.400 36.200 ;
        RECT 86.200 34.100 86.600 34.200 ;
        RECT 87.000 34.100 87.400 34.200 ;
        RECT 86.200 33.800 87.400 34.100 ;
        RECT 91.800 32.100 92.200 37.900 ;
        RECT 93.400 34.800 93.800 35.200 ;
        RECT 93.400 34.200 93.700 34.800 ;
        RECT 93.400 33.800 93.800 34.200 ;
        RECT 96.600 32.100 97.000 37.900 ;
        RECT 99.000 36.800 99.400 37.200 ;
        RECT 97.400 34.800 97.800 35.200 ;
        RECT 97.400 34.200 97.700 34.800 ;
        RECT 97.400 33.800 97.800 34.200 ;
        RECT 98.200 33.100 98.600 35.900 ;
        RECT 99.000 35.200 99.300 36.800 ;
        RECT 99.000 34.800 99.400 35.200 ;
        RECT 99.000 33.200 99.300 34.800 ;
        RECT 99.800 34.200 100.100 54.800 ;
        RECT 100.600 52.100 101.000 57.900 ;
        RECT 101.400 57.800 101.800 58.200 ;
        RECT 103.000 57.200 103.300 66.800 ;
        RECT 104.600 65.200 104.900 73.800 ;
        RECT 105.400 73.100 105.800 75.900 ;
        RECT 108.600 75.800 109.800 76.100 ;
        RECT 111.800 75.800 112.200 76.200 ;
        RECT 111.800 75.200 112.100 75.800 ;
        RECT 111.800 74.800 112.200 75.200 ;
        RECT 112.600 74.200 112.900 93.800 ;
        RECT 115.800 93.200 116.100 93.800 ;
        RECT 115.800 92.800 116.200 93.200 ;
        RECT 113.400 83.100 113.800 88.900 ;
        RECT 115.800 88.800 116.200 89.200 ;
        RECT 115.800 88.200 116.100 88.800 ;
        RECT 114.200 86.800 114.600 87.200 ;
        RECT 114.200 86.200 114.500 86.800 ;
        RECT 114.200 85.800 114.600 86.200 ;
        RECT 115.000 85.100 115.400 87.900 ;
        RECT 115.800 87.800 116.200 88.200 ;
        RECT 116.600 87.100 116.900 95.800 ;
        RECT 117.400 94.800 117.800 95.200 ;
        RECT 118.200 95.100 118.500 96.800 ;
        RECT 122.200 96.200 122.500 123.800 ;
        RECT 125.400 123.100 125.800 128.900 ;
        RECT 127.000 125.100 127.400 127.900 ;
        RECT 127.800 125.100 128.200 127.900 ;
        RECT 129.400 123.100 129.800 128.900 ;
        RECT 131.000 127.800 131.400 128.200 ;
        RECT 131.000 126.200 131.300 127.800 ;
        RECT 131.000 125.800 131.400 126.200 ;
        RECT 131.000 124.800 131.400 125.200 ;
        RECT 123.000 121.800 123.400 122.200 ;
        RECT 123.000 119.200 123.300 121.800 ;
        RECT 123.800 119.800 124.200 120.200 ;
        RECT 123.000 118.800 123.400 119.200 ;
        RECT 123.800 115.200 124.100 119.800 ;
        RECT 129.400 117.800 129.800 118.200 ;
        RECT 129.400 117.200 129.700 117.800 ;
        RECT 129.400 116.800 129.800 117.200 ;
        RECT 123.800 114.800 124.200 115.200 ;
        RECT 124.600 114.800 125.000 115.200 ;
        RECT 129.400 115.100 129.800 115.200 ;
        RECT 130.200 115.100 130.600 115.200 ;
        RECT 129.400 114.800 130.600 115.100 ;
        RECT 123.800 113.800 124.200 114.200 ;
        RECT 123.800 110.200 124.100 113.800 ;
        RECT 124.600 111.200 124.900 114.800 ;
        RECT 131.000 114.200 131.300 124.800 ;
        RECT 134.200 123.100 134.600 128.900 ;
        RECT 135.000 124.800 135.400 125.200 ;
        RECT 135.000 124.200 135.300 124.800 ;
        RECT 135.000 123.800 135.400 124.200 ;
        RECT 132.600 116.800 133.000 117.200 ;
        RECT 132.600 116.200 132.900 116.800 ;
        RECT 132.600 115.800 133.000 116.200 ;
        RECT 125.400 113.800 125.800 114.200 ;
        RECT 129.400 114.100 129.800 114.200 ;
        RECT 130.200 114.100 130.600 114.200 ;
        RECT 129.400 113.800 130.600 114.100 ;
        RECT 131.000 113.800 131.400 114.200 ;
        RECT 131.800 114.100 132.200 114.200 ;
        RECT 132.600 114.100 133.000 114.200 ;
        RECT 131.800 113.800 133.000 114.100 ;
        RECT 124.600 110.800 125.000 111.200 ;
        RECT 123.800 109.800 124.200 110.200 ;
        RECT 124.600 103.100 125.000 108.900 ;
        RECT 125.400 99.200 125.700 113.800 ;
        RECT 131.000 113.200 131.300 113.800 ;
        RECT 126.200 113.100 126.600 113.200 ;
        RECT 127.000 113.100 127.400 113.200 ;
        RECT 126.200 112.800 127.400 113.100 ;
        RECT 131.000 112.800 131.400 113.200 ;
        RECT 133.400 112.100 133.800 112.200 ;
        RECT 134.200 112.100 134.600 112.200 ;
        RECT 133.400 111.800 134.600 112.100 ;
        RECT 127.000 110.800 127.400 111.200 ;
        RECT 127.000 109.200 127.300 110.800 ;
        RECT 127.800 109.800 128.200 110.200 ;
        RECT 127.000 108.800 127.400 109.200 ;
        RECT 126.200 100.800 126.600 101.200 ;
        RECT 123.800 98.800 124.200 99.200 ;
        RECT 125.400 98.800 125.800 99.200 ;
        RECT 123.800 98.200 124.100 98.800 ;
        RECT 123.800 97.800 124.200 98.200 ;
        RECT 119.000 96.100 119.400 96.200 ;
        RECT 119.800 96.100 120.200 96.200 ;
        RECT 119.000 95.800 120.200 96.100 ;
        RECT 122.200 95.800 122.600 96.200 ;
        RECT 122.200 95.200 122.500 95.800 ;
        RECT 126.200 95.200 126.500 100.800 ;
        RECT 127.800 100.200 128.100 109.800 ;
        RECT 131.000 109.100 131.400 109.200 ;
        RECT 131.800 109.100 132.200 109.200 ;
        RECT 131.000 108.800 132.200 109.100 ;
        RECT 134.200 107.800 134.600 108.200 ;
        RECT 129.400 106.800 129.800 107.200 ;
        RECT 131.800 107.100 132.200 107.200 ;
        RECT 132.600 107.100 133.000 107.200 ;
        RECT 131.800 106.800 133.000 107.100 ;
        RECT 129.400 106.200 129.700 106.800 ;
        RECT 129.400 105.800 129.800 106.200 ;
        RECT 127.800 99.800 128.200 100.200 ;
        RECT 127.800 99.200 128.100 99.800 ;
        RECT 127.800 98.800 128.200 99.200 ;
        RECT 118.200 94.800 119.300 95.100 ;
        RECT 122.200 94.800 122.600 95.200 ;
        RECT 125.400 94.800 125.800 95.200 ;
        RECT 126.200 94.800 126.600 95.200 ;
        RECT 117.400 94.200 117.700 94.800 ;
        RECT 119.000 94.200 119.300 94.800 ;
        RECT 117.400 93.800 117.800 94.200 ;
        RECT 119.000 93.800 119.400 94.200 ;
        RECT 122.200 94.100 122.600 94.200 ;
        RECT 123.000 94.100 123.400 94.200 ;
        RECT 122.200 93.800 123.400 94.100 ;
        RECT 125.400 92.200 125.700 94.800 ;
        RECT 127.000 93.800 127.400 94.200 ;
        RECT 125.400 91.800 125.800 92.200 ;
        RECT 125.400 90.200 125.700 91.800 ;
        RECT 125.400 89.800 125.800 90.200 ;
        RECT 117.400 87.100 117.800 87.200 ;
        RECT 116.600 86.800 117.800 87.100 ;
        RECT 116.600 85.800 117.000 86.200 ;
        RECT 118.200 86.100 118.600 86.200 ;
        RECT 119.000 86.100 119.400 86.200 ;
        RECT 118.200 85.800 119.400 86.100 ;
        RECT 116.600 85.200 116.900 85.800 ;
        RECT 116.600 84.800 117.000 85.200 ;
        RECT 119.000 84.200 119.300 85.800 ;
        RECT 119.000 83.800 119.400 84.200 ;
        RECT 115.800 82.800 116.200 83.200 ;
        RECT 121.400 83.100 121.800 88.900 ;
        RECT 122.200 86.800 122.600 87.200 ;
        RECT 125.400 86.800 125.800 87.200 ;
        RECT 122.200 86.200 122.500 86.800 ;
        RECT 125.400 86.300 125.700 86.800 ;
        RECT 122.200 85.800 122.600 86.200 ;
        RECT 125.400 85.900 125.800 86.300 ;
        RECT 115.800 79.200 116.100 82.800 ;
        RECT 114.200 79.100 114.600 79.200 ;
        RECT 115.000 79.100 115.400 79.200 ;
        RECT 114.200 78.800 115.400 79.100 ;
        RECT 115.800 78.800 116.200 79.200 ;
        RECT 115.800 76.200 116.100 78.800 ;
        RECT 118.200 77.800 118.600 78.200 ;
        RECT 113.400 75.800 113.800 76.200 ;
        RECT 115.800 75.800 116.200 76.200 ;
        RECT 107.000 74.100 107.400 74.200 ;
        RECT 107.800 74.100 108.200 74.200 ;
        RECT 107.000 73.800 108.200 74.100 ;
        RECT 112.600 73.800 113.000 74.200 ;
        RECT 113.400 73.200 113.700 75.800 ;
        RECT 115.000 74.800 115.400 75.200 ;
        RECT 115.800 75.100 116.200 75.200 ;
        RECT 116.600 75.100 117.000 75.200 ;
        RECT 115.800 74.800 117.000 75.100 ;
        RECT 115.000 73.200 115.300 74.800 ;
        RECT 118.200 74.200 118.500 77.800 ;
        RECT 119.000 77.100 119.400 77.200 ;
        RECT 119.800 77.100 120.200 77.200 ;
        RECT 119.000 76.800 120.200 77.100 ;
        RECT 118.200 73.800 118.600 74.200 ;
        RECT 109.400 73.100 109.800 73.200 ;
        RECT 110.200 73.100 110.600 73.200 ;
        RECT 109.400 72.800 110.600 73.100 ;
        RECT 113.400 72.800 113.800 73.200 ;
        RECT 115.000 72.800 115.400 73.200 ;
        RECT 115.800 72.800 116.200 73.200 ;
        RECT 106.200 69.800 106.600 70.200 ;
        RECT 106.200 67.200 106.500 69.800 ;
        RECT 115.800 69.200 116.100 72.800 ;
        RECT 121.400 72.100 121.800 77.900 ;
        RECT 122.200 75.200 122.500 85.800 ;
        RECT 126.200 83.100 126.600 88.900 ;
        RECT 127.000 87.200 127.300 93.800 ;
        RECT 129.400 93.100 129.800 95.900 ;
        RECT 130.200 93.800 130.600 94.200 ;
        RECT 130.200 93.200 130.500 93.800 ;
        RECT 130.200 92.800 130.600 93.200 ;
        RECT 131.000 92.100 131.400 97.900 ;
        RECT 131.800 90.200 132.100 106.800 ;
        RECT 134.200 106.200 134.500 107.800 ;
        RECT 135.800 107.200 136.100 134.800 ;
        RECT 136.600 134.200 136.900 134.800 ;
        RECT 136.600 133.800 137.000 134.200 ;
        RECT 138.200 134.100 138.600 134.200 ;
        RECT 139.000 134.100 139.400 134.200 ;
        RECT 138.200 133.800 139.400 134.100 ;
        RECT 139.800 130.200 140.100 134.800 ;
        RECT 139.800 129.800 140.200 130.200 ;
        RECT 136.600 129.100 137.000 129.200 ;
        RECT 137.400 129.100 137.800 129.200 ;
        RECT 136.600 128.800 137.800 129.100 ;
        RECT 139.000 127.800 139.400 128.200 ;
        RECT 139.000 127.200 139.300 127.800 ;
        RECT 137.400 127.100 137.800 127.200 ;
        RECT 138.200 127.100 138.600 127.200 ;
        RECT 137.400 126.800 138.600 127.100 ;
        RECT 139.000 126.800 139.400 127.200 ;
        RECT 140.600 126.200 140.900 137.800 ;
        RECT 142.200 135.200 142.500 143.800 ;
        RECT 143.800 135.200 144.100 144.800 ;
        RECT 145.400 144.800 145.800 145.200 ;
        RECT 146.200 145.100 146.600 145.200 ;
        RECT 147.000 145.100 147.400 145.200 ;
        RECT 146.200 144.800 147.400 145.100 ;
        RECT 145.400 143.200 145.700 144.800 ;
        RECT 148.600 144.200 148.900 145.800 ;
        RECT 148.600 143.800 149.000 144.200 ;
        RECT 145.400 142.800 145.800 143.200 ;
        RECT 149.400 142.200 149.700 146.800 ;
        RECT 144.600 141.800 145.000 142.200 ;
        RECT 145.400 141.800 145.800 142.200 ;
        RECT 149.400 141.800 149.800 142.200 ;
        RECT 144.600 137.200 144.900 141.800 ;
        RECT 145.400 139.200 145.700 141.800 ;
        RECT 155.000 139.200 155.300 146.800 ;
        RECT 155.800 146.800 156.200 147.200 ;
        RECT 159.800 146.800 160.200 147.200 ;
        RECT 155.800 141.200 156.100 146.800 ;
        RECT 157.400 145.800 157.800 146.200 ;
        RECT 159.000 145.800 159.400 146.200 ;
        RECT 157.400 145.200 157.700 145.800 ;
        RECT 159.000 145.200 159.300 145.800 ;
        RECT 157.400 144.800 157.800 145.200 ;
        RECT 159.000 144.800 159.400 145.200 ;
        RECT 161.400 141.800 161.800 142.200 ;
        RECT 155.800 140.800 156.200 141.200 ;
        RECT 161.400 139.200 161.700 141.800 ;
        RECT 145.400 138.800 145.800 139.200 ;
        RECT 148.600 138.800 149.000 139.200 ;
        RECT 155.000 138.800 155.400 139.200 ;
        RECT 161.400 138.800 161.800 139.200 ;
        RECT 144.600 136.800 145.000 137.200 ;
        RECT 148.600 136.200 148.900 138.800 ;
        RECT 148.600 136.100 149.000 136.200 ;
        RECT 149.400 136.100 149.800 136.200 ;
        RECT 148.600 135.800 149.800 136.100 ;
        RECT 142.200 135.100 142.600 135.200 ;
        RECT 143.000 135.100 143.400 135.200 ;
        RECT 142.200 134.800 143.400 135.100 ;
        RECT 143.800 134.800 144.200 135.200 ;
        RECT 146.200 134.800 146.600 135.200 ;
        RECT 146.200 134.200 146.500 134.800 ;
        RECT 146.200 133.800 146.600 134.200 ;
        RECT 146.200 131.200 146.500 133.800 ;
        RECT 151.800 133.100 152.200 135.900 ;
        RECT 152.600 134.800 153.000 135.200 ;
        RECT 152.600 134.200 152.900 134.800 ;
        RECT 152.600 133.800 153.000 134.200 ;
        RECT 153.400 132.100 153.800 137.900 ;
        RECT 156.600 134.800 157.000 135.200 ;
        RECT 156.600 132.200 156.900 134.800 ;
        RECT 156.600 131.800 157.000 132.200 ;
        RECT 158.200 132.100 158.600 137.900 ;
        RECT 161.400 137.800 161.800 138.200 ;
        RECT 161.400 136.200 161.700 137.800 ;
        RECT 161.400 135.800 161.800 136.200 ;
        RECT 161.400 135.200 161.700 135.800 ;
        RECT 161.400 134.800 161.800 135.200 ;
        RECT 163.000 133.200 163.300 149.800 ;
        RECT 169.400 149.100 169.800 149.200 ;
        RECT 170.200 149.100 170.600 149.200 ;
        RECT 169.400 148.800 170.600 149.100 ;
        RECT 171.000 148.800 171.400 149.200 ;
        RECT 173.400 148.800 173.800 149.200 ;
        RECT 174.200 148.800 174.600 149.200 ;
        RECT 167.800 147.800 168.200 148.200 ;
        RECT 168.600 147.800 169.000 148.200 ;
        RECT 164.600 146.800 165.000 147.200 ;
        RECT 163.800 144.800 164.200 145.200 ;
        RECT 163.800 144.200 164.100 144.800 ;
        RECT 163.800 143.800 164.200 144.200 ;
        RECT 164.600 137.200 164.900 146.800 ;
        RECT 167.000 144.800 167.400 145.200 ;
        RECT 167.000 142.200 167.300 144.800 ;
        RECT 167.000 141.800 167.400 142.200 ;
        RECT 164.600 136.800 165.000 137.200 ;
        RECT 166.200 135.800 166.600 136.200 ;
        RECT 166.200 135.200 166.500 135.800 ;
        RECT 163.800 135.100 164.200 135.200 ;
        RECT 164.600 135.100 165.000 135.200 ;
        RECT 163.800 134.800 165.000 135.100 ;
        RECT 165.400 134.800 165.800 135.200 ;
        RECT 166.200 134.800 166.600 135.200 ;
        RECT 165.400 133.200 165.700 134.800 ;
        RECT 161.400 132.800 161.800 133.200 ;
        RECT 163.000 132.800 163.400 133.200 ;
        RECT 163.800 132.800 164.200 133.200 ;
        RECT 165.400 132.800 165.800 133.200 ;
        RECT 161.400 132.100 161.700 132.800 ;
        RECT 163.800 132.100 164.100 132.800 ;
        RECT 161.400 131.800 164.100 132.100 ;
        RECT 146.200 130.800 146.600 131.200 ;
        RECT 160.600 129.800 161.000 130.200 ;
        RECT 142.200 128.800 142.600 129.200 ;
        RECT 144.600 129.100 145.000 129.200 ;
        RECT 145.400 129.100 145.800 129.200 ;
        RECT 144.600 128.800 145.800 129.100 ;
        RECT 142.200 127.200 142.500 128.800 ;
        RECT 142.200 126.800 142.600 127.200 ;
        RECT 138.200 126.100 138.600 126.200 ;
        RECT 139.000 126.100 139.400 126.200 ;
        RECT 138.200 125.800 139.400 126.100 ;
        RECT 140.600 125.800 141.000 126.200 ;
        RECT 140.600 125.200 140.900 125.800 ;
        RECT 140.600 124.800 141.000 125.200 ;
        RECT 142.200 124.800 142.600 125.200 ;
        RECT 138.200 115.800 138.600 116.200 ;
        RECT 138.200 115.200 138.500 115.800 ;
        RECT 138.200 114.800 138.600 115.200 ;
        RECT 139.000 112.100 139.400 118.900 ;
        RECT 139.800 112.100 140.200 118.900 ;
        RECT 140.600 112.100 141.000 118.900 ;
        RECT 141.400 112.100 141.800 117.900 ;
        RECT 142.200 113.200 142.500 124.800 ;
        RECT 147.000 123.100 147.400 128.900 ;
        RECT 151.000 126.800 151.400 127.200 ;
        RECT 151.000 126.300 151.300 126.800 ;
        RECT 147.800 125.800 148.200 126.200 ;
        RECT 151.000 125.900 151.400 126.300 ;
        RECT 147.800 125.200 148.100 125.800 ;
        RECT 147.800 124.800 148.200 125.200 ;
        RECT 143.800 121.800 144.200 122.200 ;
        RECT 144.600 121.800 145.000 122.200 ;
        RECT 142.200 112.800 142.600 113.200 ;
        RECT 143.000 112.100 143.400 117.900 ;
        RECT 143.800 116.200 144.100 121.800 ;
        RECT 144.600 120.200 144.900 121.800 ;
        RECT 144.600 119.800 145.000 120.200 ;
        RECT 143.800 115.800 144.200 116.200 ;
        RECT 143.800 114.800 144.200 115.200 ;
        RECT 143.800 114.200 144.100 114.800 ;
        RECT 143.800 113.800 144.200 114.200 ;
        RECT 144.600 112.100 145.000 117.900 ;
        RECT 145.400 112.100 145.800 118.900 ;
        RECT 146.200 112.100 146.600 118.900 ;
        RECT 137.400 108.100 137.800 108.200 ;
        RECT 138.200 108.100 138.600 108.200 ;
        RECT 137.400 107.800 138.600 108.100 ;
        RECT 135.800 106.800 136.200 107.200 ;
        RECT 136.600 107.100 137.000 107.200 ;
        RECT 137.400 107.100 137.800 107.200 ;
        RECT 136.600 106.800 137.800 107.100 ;
        RECT 132.600 105.800 133.000 106.200 ;
        RECT 133.400 105.800 133.800 106.200 ;
        RECT 134.200 105.800 134.600 106.200 ;
        RECT 136.600 106.100 137.000 106.200 ;
        RECT 137.400 106.100 137.800 106.200 ;
        RECT 136.600 105.800 137.800 106.100 ;
        RECT 132.600 102.200 132.900 105.800 ;
        RECT 133.400 105.200 133.700 105.800 ;
        RECT 133.400 104.800 133.800 105.200 ;
        RECT 135.000 104.800 135.400 105.200 ;
        RECT 132.600 101.800 133.000 102.200 ;
        RECT 132.600 94.800 133.000 95.200 ;
        RECT 132.600 93.200 132.900 94.800 ;
        RECT 132.600 92.800 133.000 93.200 ;
        RECT 134.200 91.800 134.600 92.200 ;
        RECT 130.200 89.800 130.600 90.200 ;
        RECT 131.800 89.800 132.200 90.200 ;
        RECT 133.400 89.800 133.800 90.200 ;
        RECT 127.000 86.800 127.400 87.200 ;
        RECT 127.800 85.100 128.200 87.900 ;
        RECT 128.600 87.800 129.000 88.200 ;
        RECT 128.600 86.200 128.900 87.800 ;
        RECT 130.200 86.200 130.500 89.800 ;
        RECT 133.400 87.200 133.700 89.800 ;
        RECT 131.000 87.100 131.400 87.200 ;
        RECT 131.800 87.100 132.200 87.200 ;
        RECT 131.000 86.800 132.200 87.100 ;
        RECT 133.400 86.800 133.800 87.200 ;
        RECT 134.200 86.200 134.500 91.800 ;
        RECT 135.000 89.200 135.300 104.800 ;
        RECT 136.600 102.200 136.900 105.800 ;
        RECT 139.800 103.800 140.200 104.200 ;
        RECT 136.600 101.800 137.000 102.200 ;
        RECT 135.800 92.100 136.200 97.900 ;
        RECT 139.800 95.200 140.100 103.800 ;
        RECT 142.200 103.100 142.600 108.900 ;
        RECT 145.400 106.800 145.800 107.200 ;
        RECT 145.400 106.200 145.700 106.800 ;
        RECT 145.400 105.800 145.800 106.200 ;
        RECT 147.000 103.100 147.400 108.900 ;
        RECT 147.800 107.200 148.100 124.800 ;
        RECT 151.800 123.100 152.200 128.900 ;
        RECT 154.200 128.800 154.600 129.200 ;
        RECT 154.200 128.200 154.500 128.800 ;
        RECT 153.400 125.100 153.800 127.900 ;
        RECT 154.200 127.800 154.600 128.200 ;
        RECT 157.400 127.100 157.800 127.200 ;
        RECT 158.200 127.100 158.600 127.200 ;
        RECT 157.400 126.800 158.600 127.100 ;
        RECT 159.800 126.800 160.200 127.200 ;
        RECT 159.800 126.200 160.100 126.800 ;
        RECT 160.600 126.200 160.900 129.800 ;
        RECT 161.400 128.100 161.800 128.200 ;
        RECT 162.200 128.100 162.600 128.200 ;
        RECT 161.400 127.800 162.600 128.100 ;
        RECT 164.600 127.800 165.000 128.200 ;
        RECT 164.600 127.200 164.900 127.800 ;
        RECT 161.400 127.100 161.800 127.200 ;
        RECT 162.200 127.100 162.600 127.200 ;
        RECT 161.400 126.800 162.600 127.100 ;
        RECT 163.000 126.800 163.400 127.200 ;
        RECT 164.600 126.800 165.000 127.200 ;
        RECT 157.400 126.100 157.800 126.200 ;
        RECT 158.200 126.100 158.600 126.200 ;
        RECT 157.400 125.800 158.600 126.100 ;
        RECT 159.800 125.800 160.200 126.200 ;
        RECT 160.600 125.800 161.000 126.200 ;
        RECT 162.200 125.800 162.600 126.200 ;
        RECT 159.800 121.200 160.100 125.800 ;
        RECT 159.800 120.800 160.200 121.200 ;
        RECT 149.400 117.800 149.800 118.200 ;
        RECT 149.400 115.200 149.700 117.800 ;
        RECT 162.200 117.200 162.500 125.800 ;
        RECT 163.000 123.200 163.300 126.800 ;
        RECT 166.200 126.200 166.500 134.800 ;
        RECT 167.800 134.200 168.100 147.800 ;
        RECT 168.600 147.200 168.900 147.800 ;
        RECT 171.000 147.200 171.300 148.800 ;
        RECT 173.400 147.200 173.700 148.800 ;
        RECT 174.200 148.200 174.500 148.800 ;
        RECT 174.200 147.800 174.600 148.200 ;
        RECT 168.600 146.800 169.000 147.200 ;
        RECT 171.000 146.800 171.400 147.200 ;
        RECT 171.800 146.800 172.200 147.200 ;
        RECT 173.400 146.800 173.800 147.200 ;
        RECT 171.000 145.800 171.400 146.200 ;
        RECT 171.000 142.200 171.300 145.800 ;
        RECT 171.800 145.200 172.100 146.800 ;
        RECT 176.600 146.200 176.900 151.800 ;
        RECT 177.400 151.200 177.700 151.800 ;
        RECT 177.400 150.800 177.800 151.200 ;
        RECT 178.200 150.200 178.500 154.800 ;
        RECT 180.600 153.200 180.900 154.800 ;
        RECT 179.000 152.800 179.400 153.200 ;
        RECT 179.800 153.100 180.200 153.200 ;
        RECT 180.600 153.100 181.000 153.200 ;
        RECT 179.800 152.800 181.000 153.100 ;
        RECT 178.200 149.800 178.600 150.200 ;
        RECT 177.400 147.800 177.800 148.200 ;
        RECT 177.400 147.200 177.700 147.800 ;
        RECT 177.400 146.800 177.800 147.200 ;
        RECT 176.600 145.800 177.000 146.200 ;
        RECT 171.800 144.800 172.200 145.200 ;
        RECT 173.400 144.800 173.800 145.200 ;
        RECT 171.000 141.800 171.400 142.200 ;
        RECT 172.600 141.800 173.000 142.200 ;
        RECT 172.600 141.200 172.900 141.800 ;
        RECT 171.800 140.800 172.200 141.200 ;
        RECT 172.600 140.800 173.000 141.200 ;
        RECT 170.200 137.800 170.600 138.200 ;
        RECT 170.200 136.200 170.500 137.800 ;
        RECT 170.200 135.800 170.600 136.200 ;
        RECT 171.800 135.200 172.100 140.800 ;
        RECT 172.600 140.100 173.000 140.200 ;
        RECT 173.400 140.100 173.700 144.800 ;
        RECT 172.600 139.800 173.700 140.100 ;
        RECT 175.000 142.800 175.400 143.200 ;
        RECT 172.600 137.800 173.000 138.200 ;
        RECT 172.600 136.200 172.900 137.800 ;
        RECT 175.000 137.200 175.300 142.800 ;
        RECT 176.600 141.200 176.900 145.800 ;
        RECT 178.200 143.100 178.500 149.800 ;
        RECT 179.000 146.200 179.300 152.800 ;
        RECT 181.400 149.200 181.700 161.800 ;
        RECT 184.600 156.800 185.000 157.200 ;
        RECT 184.600 156.200 184.900 156.800 ;
        RECT 184.600 155.800 185.000 156.200 ;
        RECT 188.600 155.200 188.900 165.800 ;
        RECT 192.700 165.100 193.000 167.500 ;
        RECT 193.400 167.400 193.800 167.500 ;
        RECT 195.100 167.400 195.500 167.500 ;
        RECT 195.900 167.100 196.200 167.500 ;
        RECT 198.200 167.800 198.600 168.200 ;
        RECT 193.400 166.800 196.200 167.100 ;
        RECT 193.400 166.100 193.700 166.800 ;
        RECT 193.300 165.700 193.700 166.100 ;
        RECT 195.900 165.100 196.200 166.800 ;
        RECT 192.700 164.700 193.100 165.100 ;
        RECT 195.800 164.700 196.200 165.100 ;
        RECT 196.600 166.800 197.000 167.200 ;
        RECT 197.400 166.800 197.800 167.200 ;
        RECT 196.600 164.200 196.900 166.800 ;
        RECT 197.400 165.200 197.700 166.800 ;
        RECT 198.200 166.200 198.500 167.800 ;
        RECT 198.200 165.800 198.600 166.200 ;
        RECT 199.000 166.100 199.400 166.200 ;
        RECT 199.800 166.100 200.200 166.200 ;
        RECT 199.000 165.800 200.200 166.100 ;
        RECT 201.400 165.800 201.800 166.200 ;
        RECT 201.400 165.200 201.700 165.800 ;
        RECT 197.400 164.800 197.800 165.200 ;
        RECT 199.800 164.800 200.200 165.200 ;
        RECT 201.400 164.800 201.800 165.200 ;
        RECT 196.600 163.800 197.000 164.200 ;
        RECT 195.800 157.800 196.200 158.200 ;
        RECT 190.200 155.800 190.600 156.200 ;
        RECT 190.200 155.200 190.500 155.800 ;
        RECT 184.600 154.800 185.000 155.200 ;
        RECT 188.600 154.800 189.000 155.200 ;
        RECT 189.400 154.800 189.800 155.200 ;
        RECT 190.200 154.800 190.600 155.200 ;
        RECT 183.000 154.100 183.400 154.200 ;
        RECT 183.800 154.100 184.200 154.200 ;
        RECT 183.000 153.800 184.200 154.100 ;
        RECT 183.000 152.800 183.400 153.200 ;
        RECT 182.200 151.800 182.600 152.200 ;
        RECT 181.400 148.800 181.800 149.200 ;
        RECT 182.200 149.100 182.500 151.800 ;
        RECT 183.000 150.200 183.300 152.800 ;
        RECT 183.800 151.800 184.200 152.200 ;
        RECT 183.000 149.800 183.400 150.200 ;
        RECT 183.800 149.200 184.100 151.800 ;
        RECT 184.600 151.200 184.900 154.800 ;
        RECT 189.400 154.200 189.700 154.800 ;
        RECT 188.600 153.800 189.000 154.200 ;
        RECT 189.400 153.800 189.800 154.200 ;
        RECT 194.200 153.800 194.600 154.200 ;
        RECT 188.600 153.100 188.900 153.800 ;
        RECT 188.600 152.800 189.700 153.100 ;
        RECT 187.800 151.800 188.200 152.200 ;
        RECT 184.600 150.800 185.000 151.200 ;
        RECT 182.200 148.800 183.300 149.100 ;
        RECT 183.800 148.800 184.200 149.200 ;
        RECT 183.000 148.200 183.300 148.800 ;
        RECT 187.800 148.200 188.100 151.800 ;
        RECT 189.400 149.200 189.700 152.800 ;
        RECT 191.800 151.800 192.200 152.200 ;
        RECT 191.800 150.200 192.100 151.800 ;
        RECT 194.200 151.200 194.500 153.800 ;
        RECT 195.000 153.100 195.400 155.900 ;
        RECT 195.800 154.200 196.100 157.800 ;
        RECT 195.800 153.800 196.200 154.200 ;
        RECT 196.600 152.100 197.000 157.900 ;
        RECT 198.200 154.800 198.600 155.200 ;
        RECT 194.200 150.800 194.600 151.200 ;
        RECT 196.600 150.800 197.000 151.200 ;
        RECT 191.800 149.800 192.200 150.200 ;
        RECT 196.600 149.200 196.900 150.800 ;
        RECT 189.400 148.800 189.800 149.200 ;
        RECT 191.000 148.800 191.400 149.200 ;
        RECT 196.600 148.800 197.000 149.200 ;
        RECT 191.000 148.200 191.300 148.800 ;
        RECT 181.400 147.800 181.800 148.200 ;
        RECT 182.200 147.800 182.600 148.200 ;
        RECT 183.000 147.800 183.400 148.200 ;
        RECT 184.600 147.800 185.000 148.200 ;
        RECT 187.800 147.800 188.200 148.200 ;
        RECT 191.000 147.800 191.400 148.200 ;
        RECT 195.000 148.100 195.400 148.200 ;
        RECT 195.800 148.100 196.200 148.200 ;
        RECT 195.000 147.800 196.200 148.100 ;
        RECT 179.000 145.800 179.400 146.200 ;
        RECT 179.800 145.800 180.200 146.200 ;
        RECT 179.000 145.200 179.300 145.800 ;
        RECT 179.000 144.800 179.400 145.200 ;
        RECT 177.400 142.800 178.500 143.100 ;
        RECT 176.600 140.800 177.000 141.200 ;
        RECT 175.800 138.800 176.200 139.200 ;
        RECT 175.800 138.200 176.100 138.800 ;
        RECT 175.800 137.800 176.200 138.200 ;
        RECT 175.000 136.800 175.400 137.200 ;
        RECT 176.600 136.800 177.000 137.200 ;
        RECT 172.600 135.800 173.000 136.200 ;
        RECT 168.600 134.800 169.000 135.200 ;
        RECT 171.800 134.800 172.200 135.200 ;
        RECT 173.400 135.100 173.800 135.200 ;
        RECT 174.200 135.100 174.600 135.200 ;
        RECT 173.400 134.800 174.600 135.100 ;
        RECT 167.800 133.800 168.200 134.200 ;
        RECT 167.000 132.100 167.400 132.200 ;
        RECT 167.800 132.100 168.200 132.200 ;
        RECT 167.000 131.800 168.200 132.100 ;
        RECT 168.600 130.200 168.900 134.800 ;
        RECT 175.000 134.200 175.300 136.800 ;
        RECT 175.000 133.800 175.400 134.200 ;
        RECT 176.600 132.200 176.900 136.800 ;
        RECT 177.400 135.200 177.700 142.800 ;
        RECT 178.200 141.800 178.600 142.200 ;
        RECT 178.200 137.200 178.500 141.800 ;
        RECT 178.200 136.800 178.600 137.200 ;
        RECT 178.200 136.100 178.600 136.200 ;
        RECT 179.000 136.100 179.400 136.200 ;
        RECT 178.200 135.800 179.400 136.100 ;
        RECT 179.800 135.200 180.100 145.800 ;
        RECT 180.600 144.800 181.000 145.200 ;
        RECT 180.600 144.200 180.900 144.800 ;
        RECT 180.600 143.800 181.000 144.200 ;
        RECT 180.600 135.800 181.000 136.200 ;
        RECT 180.600 135.200 180.900 135.800 ;
        RECT 177.400 134.800 177.800 135.200 ;
        RECT 178.200 135.100 178.600 135.200 ;
        RECT 179.000 135.100 179.400 135.200 ;
        RECT 178.200 134.800 179.400 135.100 ;
        RECT 179.800 134.800 180.200 135.200 ;
        RECT 180.600 134.800 181.000 135.200 ;
        RECT 178.200 134.100 178.600 134.200 ;
        RECT 179.000 134.100 179.400 134.200 ;
        RECT 178.200 133.800 179.400 134.100 ;
        RECT 179.800 134.100 180.200 134.200 ;
        RECT 180.600 134.100 181.000 134.200 ;
        RECT 179.800 133.800 181.000 134.100 ;
        RECT 181.400 133.200 181.700 147.800 ;
        RECT 182.200 147.200 182.500 147.800 ;
        RECT 184.600 147.200 184.900 147.800 ;
        RECT 182.200 146.800 182.600 147.200 ;
        RECT 183.000 146.800 183.400 147.200 ;
        RECT 184.600 146.800 185.000 147.200 ;
        RECT 187.800 147.100 188.200 147.200 ;
        RECT 188.600 147.100 189.000 147.200 ;
        RECT 187.800 146.800 189.000 147.100 ;
        RECT 182.200 145.800 182.600 146.200 ;
        RECT 182.200 145.200 182.500 145.800 ;
        RECT 182.200 144.800 182.600 145.200 ;
        RECT 183.000 140.200 183.300 146.800 ;
        RECT 185.400 145.800 185.800 146.200 ;
        RECT 186.200 146.100 186.600 146.200 ;
        RECT 187.000 146.100 187.400 146.200 ;
        RECT 186.200 145.800 187.400 146.100 ;
        RECT 187.800 146.100 188.200 146.200 ;
        RECT 188.600 146.100 189.000 146.200 ;
        RECT 187.800 145.800 189.000 146.100 ;
        RECT 183.000 139.800 183.400 140.200 ;
        RECT 184.600 136.800 185.000 137.200 ;
        RECT 184.600 136.200 184.900 136.800 ;
        RECT 184.600 135.800 185.000 136.200 ;
        RECT 185.400 135.200 185.700 145.800 ;
        RECT 186.200 144.100 186.600 144.200 ;
        RECT 187.000 144.100 187.400 144.200 ;
        RECT 186.200 143.800 187.400 144.100 ;
        RECT 191.000 143.200 191.300 147.800 ;
        RECT 194.200 146.800 194.600 147.200 ;
        RECT 197.400 146.800 197.800 147.200 ;
        RECT 194.200 146.200 194.500 146.800 ;
        RECT 197.400 146.200 197.700 146.800 ;
        RECT 192.600 145.800 193.000 146.200 ;
        RECT 194.200 145.800 194.600 146.200 ;
        RECT 197.400 145.800 197.800 146.200 ;
        RECT 191.000 142.800 191.400 143.200 ;
        RECT 192.600 142.200 192.900 145.800 ;
        RECT 193.400 144.800 193.800 145.200 ;
        RECT 193.400 144.200 193.700 144.800 ;
        RECT 193.400 143.800 193.800 144.200 ;
        RECT 194.200 144.100 194.600 144.200 ;
        RECT 195.000 144.100 195.400 144.200 ;
        RECT 194.200 143.800 195.400 144.100 ;
        RECT 196.600 144.100 197.000 144.200 ;
        RECT 197.400 144.100 197.800 144.200 ;
        RECT 196.600 143.800 197.800 144.100 ;
        RECT 195.000 142.800 195.400 143.200 ;
        RECT 191.000 141.800 191.400 142.200 ;
        RECT 192.600 141.800 193.000 142.200 ;
        RECT 191.000 139.200 191.300 141.800 ;
        RECT 192.600 139.800 193.000 140.200 ;
        RECT 192.600 139.200 192.900 139.800 ;
        RECT 191.000 138.800 191.400 139.200 ;
        RECT 192.600 138.800 193.000 139.200 ;
        RECT 193.400 136.800 193.800 137.200 ;
        RECT 193.400 136.200 193.700 136.800 ;
        RECT 195.000 136.200 195.300 142.800 ;
        RECT 195.800 141.800 196.200 142.200 ;
        RECT 195.800 136.200 196.100 141.800 ;
        RECT 198.200 136.200 198.500 154.800 ;
        RECT 199.800 149.200 200.100 164.800 ;
        RECT 202.200 164.200 202.500 172.800 ;
        RECT 203.800 168.800 204.200 169.200 ;
        RECT 203.800 168.200 204.100 168.800 ;
        RECT 203.800 167.800 204.200 168.200 ;
        RECT 204.600 167.800 205.000 168.200 ;
        RECT 204.600 167.200 204.900 167.800 ;
        RECT 204.600 166.800 205.000 167.200 ;
        RECT 202.200 163.800 202.600 164.200 ;
        RECT 201.400 152.100 201.800 157.900 ;
        RECT 199.800 148.800 200.200 149.200 ;
        RECT 202.200 148.200 202.500 163.800 ;
        RECT 203.800 151.800 204.200 152.200 ;
        RECT 202.200 147.800 202.600 148.200 ;
        RECT 202.200 147.200 202.500 147.800 ;
        RECT 202.200 146.800 202.600 147.200 ;
        RECT 199.000 144.800 199.400 145.200 ;
        RECT 199.000 143.200 199.300 144.800 ;
        RECT 201.400 143.800 201.800 144.200 ;
        RECT 199.000 142.800 199.400 143.200 ;
        RECT 199.800 141.800 200.200 142.200 ;
        RECT 199.800 138.200 200.100 141.800 ;
        RECT 201.400 139.200 201.700 143.800 ;
        RECT 201.400 138.800 201.800 139.200 ;
        RECT 203.800 138.200 204.100 151.800 ;
        RECT 204.600 146.200 204.900 166.800 ;
        RECT 204.600 145.800 205.000 146.200 ;
        RECT 199.800 137.800 200.200 138.200 ;
        RECT 203.800 137.800 204.200 138.200 ;
        RECT 187.800 135.800 188.200 136.200 ;
        RECT 189.400 136.100 189.800 136.200 ;
        RECT 190.200 136.100 190.600 136.200 ;
        RECT 189.400 135.800 190.600 136.100 ;
        RECT 193.400 135.800 193.800 136.200 ;
        RECT 195.000 135.800 195.400 136.200 ;
        RECT 195.800 135.800 196.200 136.200 ;
        RECT 197.400 135.800 197.800 136.200 ;
        RECT 198.200 135.800 198.600 136.200 ;
        RECT 199.800 135.900 200.200 136.300 ;
        RECT 203.100 135.900 203.500 136.300 ;
        RECT 183.000 135.100 183.400 135.200 ;
        RECT 183.800 135.100 184.200 135.200 ;
        RECT 183.000 134.800 184.200 135.100 ;
        RECT 185.400 134.800 185.800 135.200 ;
        RECT 186.200 134.800 186.600 135.200 ;
        RECT 186.200 134.200 186.500 134.800 ;
        RECT 183.800 133.800 184.200 134.200 ;
        RECT 186.200 133.800 186.600 134.200 ;
        RECT 183.800 133.200 184.100 133.800 ;
        RECT 181.400 132.800 181.800 133.200 ;
        RECT 183.800 132.800 184.200 133.200 ;
        RECT 186.200 132.200 186.500 133.800 ;
        RECT 170.200 131.800 170.600 132.200 ;
        RECT 176.600 131.800 177.000 132.200 ;
        RECT 179.800 131.800 180.200 132.200 ;
        RECT 186.200 131.800 186.600 132.200 ;
        RECT 168.600 129.800 169.000 130.200 ;
        RECT 169.400 128.800 169.800 129.200 ;
        RECT 169.400 128.200 169.700 128.800 ;
        RECT 169.400 127.800 169.800 128.200 ;
        RECT 168.600 127.100 169.000 127.200 ;
        RECT 169.400 127.100 169.800 127.200 ;
        RECT 168.600 126.800 169.800 127.100 ;
        RECT 163.800 125.800 164.200 126.200 ;
        RECT 166.200 125.800 166.600 126.200 ;
        RECT 167.000 126.100 167.400 126.200 ;
        RECT 167.800 126.100 168.200 126.200 ;
        RECT 167.000 125.800 168.200 126.100 ;
        RECT 163.000 122.800 163.400 123.200 ;
        RECT 163.000 120.800 163.400 121.200 ;
        RECT 163.000 119.200 163.300 120.800 ;
        RECT 163.000 118.800 163.400 119.200 ;
        RECT 151.800 116.800 152.200 117.200 ;
        RECT 162.200 116.800 162.600 117.200 ;
        RECT 151.800 116.200 152.100 116.800 ;
        RECT 151.800 115.800 152.200 116.200 ;
        RECT 159.800 115.800 160.200 116.200 ;
        RECT 149.400 114.800 149.800 115.200 ;
        RECT 151.000 114.800 151.400 115.200 ;
        RECT 156.600 115.100 157.000 115.200 ;
        RECT 157.400 115.100 157.800 115.200 ;
        RECT 156.600 114.800 157.800 115.100 ;
        RECT 151.000 111.100 151.300 114.800 ;
        RECT 159.800 114.200 160.100 115.800 ;
        RECT 160.600 114.800 161.000 115.200 ;
        RECT 160.600 114.200 160.900 114.800 ;
        RECT 162.200 114.200 162.500 116.800 ;
        RECT 163.800 116.200 164.100 125.800 ;
        RECT 164.600 125.100 165.000 125.200 ;
        RECT 165.400 125.100 165.800 125.200 ;
        RECT 164.600 124.800 165.800 125.100 ;
        RECT 165.400 123.800 165.800 124.200 ;
        RECT 165.400 119.200 165.700 123.800 ;
        RECT 170.200 119.200 170.500 131.800 ;
        RECT 171.000 130.800 171.400 131.200 ;
        RECT 171.000 128.200 171.300 130.800 ;
        RECT 176.600 129.100 177.000 129.200 ;
        RECT 177.400 129.100 177.800 129.200 ;
        RECT 176.600 128.800 177.800 129.100 ;
        RECT 179.800 128.200 180.100 131.800 ;
        RECT 187.000 129.800 187.400 130.200 ;
        RECT 183.800 128.800 184.200 129.200 ;
        RECT 183.800 128.200 184.100 128.800 ;
        RECT 171.000 127.800 171.400 128.200 ;
        RECT 174.200 127.800 174.600 128.200 ;
        RECT 177.400 127.800 177.800 128.200 ;
        RECT 179.800 127.800 180.200 128.200 ;
        RECT 183.800 127.800 184.200 128.200 ;
        RECT 172.600 126.800 173.000 127.200 ;
        RECT 173.400 126.800 173.800 127.200 ;
        RECT 172.600 126.200 172.900 126.800 ;
        RECT 173.400 126.200 173.700 126.800 ;
        RECT 174.200 126.200 174.500 127.800 ;
        RECT 172.600 125.800 173.000 126.200 ;
        RECT 173.400 125.800 173.800 126.200 ;
        RECT 174.200 125.800 174.600 126.200 ;
        RECT 174.200 125.200 174.500 125.800 ;
        RECT 177.400 125.200 177.700 127.800 ;
        RECT 179.800 125.200 180.100 127.800 ;
        RECT 187.000 127.200 187.300 129.800 ;
        RECT 187.800 129.200 188.100 135.800 ;
        RECT 194.200 134.800 194.600 135.200 ;
        RECT 194.200 134.200 194.500 134.800 ;
        RECT 189.400 133.800 189.800 134.200 ;
        RECT 191.800 134.100 192.200 134.200 ;
        RECT 192.600 134.100 193.000 134.200 ;
        RECT 191.800 133.800 193.000 134.100 ;
        RECT 194.200 133.800 194.600 134.200 ;
        RECT 189.400 130.200 189.700 133.800 ;
        RECT 195.000 130.200 195.300 135.800 ;
        RECT 197.400 134.200 197.700 135.800 ;
        RECT 199.800 134.200 200.100 135.900 ;
        RECT 201.800 134.200 202.200 134.300 ;
        RECT 195.800 134.100 196.200 134.200 ;
        RECT 196.600 134.100 197.000 134.200 ;
        RECT 195.800 133.800 197.000 134.100 ;
        RECT 197.400 133.800 197.800 134.200 ;
        RECT 198.200 134.100 198.600 134.200 ;
        RECT 199.000 134.100 199.400 134.200 ;
        RECT 198.200 133.800 199.400 134.100 ;
        RECT 199.800 133.900 202.200 134.200 ;
        RECT 199.800 133.500 200.100 133.900 ;
        RECT 200.500 133.500 200.900 133.600 ;
        RECT 202.200 133.500 202.600 133.600 ;
        RECT 203.200 133.500 203.500 135.900 ;
        RECT 204.600 134.200 204.900 145.800 ;
        RECT 204.600 133.800 205.000 134.200 ;
        RECT 195.800 132.800 196.200 133.200 ;
        RECT 199.800 133.100 200.200 133.500 ;
        RECT 200.500 133.200 202.600 133.500 ;
        RECT 200.600 132.800 201.000 133.200 ;
        RECT 203.100 133.100 203.500 133.500 ;
        RECT 195.800 132.200 196.100 132.800 ;
        RECT 195.800 131.800 196.200 132.200 ;
        RECT 189.400 129.800 189.800 130.200 ;
        RECT 195.000 129.800 195.400 130.200 ;
        RECT 199.000 129.800 199.400 130.200 ;
        RECT 199.800 129.800 200.200 130.200 ;
        RECT 203.000 129.800 203.400 130.200 ;
        RECT 199.000 129.200 199.300 129.800 ;
        RECT 187.800 128.800 188.200 129.200 ;
        RECT 199.000 128.800 199.400 129.200 ;
        RECT 199.800 128.200 200.100 129.800 ;
        RECT 203.000 129.200 203.300 129.800 ;
        RECT 203.000 128.800 203.400 129.200 ;
        RECT 193.400 127.800 193.800 128.200 ;
        RECT 199.800 127.800 200.200 128.200 ;
        RECT 201.400 127.800 201.800 128.200 ;
        RECT 202.200 128.100 202.600 128.200 ;
        RECT 203.000 128.100 203.400 128.200 ;
        RECT 202.200 127.800 203.400 128.100 ;
        RECT 187.000 127.100 187.400 127.200 ;
        RECT 187.800 127.100 188.200 127.200 ;
        RECT 187.000 126.800 188.200 127.100 ;
        RECT 193.400 126.200 193.700 127.800 ;
        RECT 201.400 127.200 201.700 127.800 ;
        RECT 195.800 126.800 196.200 127.200 ;
        RECT 197.400 126.800 197.800 127.200 ;
        RECT 198.200 126.800 198.600 127.200 ;
        RECT 201.400 126.800 201.800 127.200 ;
        RECT 203.800 126.800 204.200 127.200 ;
        RECT 195.800 126.200 196.100 126.800 ;
        RECT 182.200 125.800 182.600 126.200 ;
        RECT 191.800 125.800 192.200 126.200 ;
        RECT 193.400 126.100 193.800 126.200 ;
        RECT 194.200 126.100 194.600 126.200 ;
        RECT 193.400 125.800 194.600 126.100 ;
        RECT 195.800 125.800 196.200 126.200 ;
        RECT 182.200 125.200 182.500 125.800 ;
        RECT 171.000 125.100 171.400 125.200 ;
        RECT 171.800 125.100 172.200 125.200 ;
        RECT 171.000 124.800 172.200 125.100 ;
        RECT 174.200 124.800 174.600 125.200 ;
        RECT 177.400 124.800 177.800 125.200 ;
        RECT 179.800 124.800 180.200 125.200 ;
        RECT 182.200 124.800 182.600 125.200 ;
        RECT 174.200 123.800 174.600 124.200 ;
        RECT 165.400 118.800 165.800 119.200 ;
        RECT 170.200 118.800 170.600 119.200 ;
        RECT 167.000 117.800 167.400 118.200 ;
        RECT 167.000 116.200 167.300 117.800 ;
        RECT 169.400 116.800 169.800 117.200 ;
        RECT 163.000 115.800 163.400 116.200 ;
        RECT 163.800 116.100 164.200 116.200 ;
        RECT 164.600 116.100 165.000 116.200 ;
        RECT 163.800 115.800 165.000 116.100 ;
        RECT 166.200 115.800 166.600 116.200 ;
        RECT 167.000 115.800 167.400 116.200 ;
        RECT 163.000 115.200 163.300 115.800 ;
        RECT 163.000 114.800 163.400 115.200 ;
        RECT 164.600 114.800 165.000 115.200 ;
        RECT 165.400 114.800 165.800 115.200 ;
        RECT 164.600 114.200 164.900 114.800 ;
        RECT 156.600 114.100 157.000 114.200 ;
        RECT 157.400 114.100 157.800 114.200 ;
        RECT 156.600 113.800 157.800 114.100 ;
        RECT 159.800 113.800 160.200 114.200 ;
        RECT 160.600 113.800 161.000 114.200 ;
        RECT 162.200 113.800 162.600 114.200 ;
        RECT 164.600 113.800 165.000 114.200 ;
        RECT 165.400 113.200 165.700 114.800 ;
        RECT 152.600 113.100 153.000 113.200 ;
        RECT 150.200 110.800 151.300 111.100 ;
        RECT 151.800 112.800 153.000 113.100 ;
        RECT 154.200 112.800 154.600 113.200 ;
        RECT 155.800 112.800 156.200 113.200 ;
        RECT 158.200 112.800 158.600 113.200 ;
        RECT 159.000 112.800 159.400 113.200 ;
        RECT 165.400 112.800 165.800 113.200 ;
        RECT 147.800 106.800 148.200 107.200 ;
        RECT 148.600 105.100 149.000 107.900 ;
        RECT 150.200 99.200 150.500 110.800 ;
        RECT 151.000 105.100 151.400 107.900 ;
        RECT 144.600 98.800 145.000 99.200 ;
        RECT 148.600 98.800 149.000 99.200 ;
        RECT 150.200 98.800 150.600 99.200 ;
        RECT 138.200 95.100 138.600 95.200 ;
        RECT 139.000 95.100 139.400 95.200 ;
        RECT 138.200 94.800 139.400 95.100 ;
        RECT 139.800 94.800 140.200 95.200 ;
        RECT 141.400 95.100 141.800 95.200 ;
        RECT 142.200 95.100 142.600 95.200 ;
        RECT 141.400 94.800 142.600 95.100 ;
        RECT 139.800 94.200 140.100 94.800 ;
        RECT 138.200 93.800 138.600 94.200 ;
        RECT 139.800 93.800 140.200 94.200 ;
        RECT 138.200 92.200 138.500 93.800 ;
        RECT 140.600 92.800 141.000 93.200 ;
        RECT 140.600 92.200 140.900 92.800 ;
        RECT 138.200 91.800 138.600 92.200 ;
        RECT 140.600 91.800 141.000 92.200 ;
        RECT 137.400 90.800 137.800 91.200 ;
        RECT 137.400 89.200 137.700 90.800 ;
        RECT 135.000 88.800 135.400 89.200 ;
        RECT 137.400 88.800 137.800 89.200 ;
        RECT 128.600 85.800 129.000 86.200 ;
        RECT 130.200 85.800 130.600 86.200 ;
        RECT 133.400 85.800 133.800 86.200 ;
        RECT 134.200 85.800 134.600 86.200 ;
        RECT 122.200 74.800 122.600 75.200 ;
        RECT 124.600 75.000 125.000 75.100 ;
        RECT 125.400 75.000 125.800 75.100 ;
        RECT 124.600 74.700 125.800 75.000 ;
        RECT 124.600 73.800 125.000 74.200 ;
        RECT 106.200 66.800 106.600 67.200 ;
        RECT 105.400 65.800 105.800 66.200 ;
        RECT 103.800 64.800 104.200 65.200 ;
        RECT 104.600 64.800 105.000 65.200 ;
        RECT 103.800 63.200 104.100 64.800 ;
        RECT 103.800 62.800 104.200 63.200 ;
        RECT 103.000 56.800 103.400 57.200 ;
        RECT 103.800 53.200 104.100 62.800 ;
        RECT 104.600 55.800 105.000 56.200 ;
        RECT 103.000 52.800 103.400 53.200 ;
        RECT 103.800 52.800 104.200 53.200 ;
        RECT 103.000 52.200 103.300 52.800 ;
        RECT 103.000 51.800 103.400 52.200 ;
        RECT 103.800 47.200 104.100 52.800 ;
        RECT 104.600 49.200 104.900 55.800 ;
        RECT 105.400 52.200 105.700 65.800 ;
        RECT 107.000 65.100 107.400 67.900 ;
        RECT 108.600 63.100 109.000 68.900 ;
        RECT 110.200 66.100 110.600 66.200 ;
        RECT 111.000 66.100 111.400 66.200 ;
        RECT 110.200 65.800 111.400 66.100 ;
        RECT 112.600 65.800 113.000 66.200 ;
        RECT 112.600 65.200 112.900 65.800 ;
        RECT 112.600 64.800 113.000 65.200 ;
        RECT 113.400 63.100 113.800 68.900 ;
        RECT 115.800 68.800 116.200 69.200 ;
        RECT 118.200 68.800 118.600 69.200 ;
        RECT 118.200 68.200 118.500 68.800 ;
        RECT 118.200 67.800 118.600 68.200 ;
        RECT 119.000 68.100 119.400 68.200 ;
        RECT 119.800 68.100 120.200 68.200 ;
        RECT 119.000 67.800 120.200 68.100 ;
        RECT 117.400 67.100 117.800 67.200 ;
        RECT 119.000 67.100 119.400 67.200 ;
        RECT 117.400 66.800 119.400 67.100 ;
        RECT 116.600 65.800 117.000 66.200 ;
        RECT 107.000 61.800 107.400 62.200 ;
        RECT 107.000 59.200 107.300 61.800 ;
        RECT 115.000 60.800 115.400 61.200 ;
        RECT 107.000 58.800 107.400 59.200 ;
        RECT 110.200 55.800 110.600 56.200 ;
        RECT 111.800 55.800 112.200 56.200 ;
        RECT 110.200 54.200 110.500 55.800 ;
        RECT 111.800 55.200 112.100 55.800 ;
        RECT 111.800 54.800 112.200 55.200 ;
        RECT 113.400 55.100 113.800 55.200 ;
        RECT 114.200 55.100 114.600 55.200 ;
        RECT 113.400 54.800 114.600 55.100 ;
        RECT 115.000 54.200 115.300 60.800 ;
        RECT 116.600 58.200 116.900 65.800 ;
        RECT 122.200 63.100 122.600 68.900 ;
        RECT 123.000 67.800 123.400 68.200 ;
        RECT 123.000 67.200 123.300 67.800 ;
        RECT 123.000 66.800 123.400 67.200 ;
        RECT 124.600 65.200 124.900 73.800 ;
        RECT 126.200 72.100 126.600 77.900 ;
        RECT 127.800 73.100 128.200 75.900 ;
        RECT 130.200 75.200 130.500 85.800 ;
        RECT 133.400 83.200 133.700 85.800 ;
        RECT 133.400 82.800 133.800 83.200 ;
        RECT 131.000 76.800 131.400 77.200 ;
        RECT 130.200 74.800 130.600 75.200 ;
        RECT 128.600 73.800 129.000 74.200 ;
        RECT 128.600 73.200 128.900 73.800 ;
        RECT 128.600 72.800 129.000 73.200 ;
        RECT 129.400 71.800 129.800 72.200 ;
        RECT 126.200 66.800 126.600 67.200 ;
        RECT 126.200 66.300 126.500 66.800 ;
        RECT 126.200 65.900 126.600 66.300 ;
        RECT 126.200 65.800 126.500 65.900 ;
        RECT 124.600 64.800 125.000 65.200 ;
        RECT 116.600 57.800 117.000 58.200 ;
        RECT 119.000 56.800 119.400 57.200 ;
        RECT 119.000 56.200 119.300 56.800 ;
        RECT 119.000 55.800 119.400 56.200 ;
        RECT 115.800 55.100 116.200 55.200 ;
        RECT 116.600 55.100 117.000 55.200 ;
        RECT 115.800 54.800 117.000 55.100 ;
        RECT 107.800 53.800 108.200 54.200 ;
        RECT 110.200 53.800 110.600 54.200 ;
        RECT 115.000 53.800 115.400 54.200 ;
        RECT 115.800 54.100 116.200 54.200 ;
        RECT 116.600 54.100 117.000 54.200 ;
        RECT 115.800 53.800 117.000 54.100 ;
        RECT 107.800 53.200 108.100 53.800 ;
        RECT 107.800 52.800 108.200 53.200 ;
        RECT 112.600 52.800 113.000 53.200 ;
        RECT 112.600 52.200 112.900 52.800 ;
        RECT 105.400 51.800 105.800 52.200 ;
        RECT 110.200 51.800 110.600 52.200 ;
        RECT 112.600 51.800 113.000 52.200 ;
        RECT 107.800 49.800 108.200 50.200 ;
        RECT 108.600 49.800 109.000 50.200 ;
        RECT 107.800 49.200 108.100 49.800 ;
        RECT 104.600 48.800 105.000 49.200 ;
        RECT 107.800 48.800 108.200 49.200 ;
        RECT 108.600 48.200 108.900 49.800 ;
        RECT 110.200 49.200 110.500 51.800 ;
        RECT 115.000 50.800 115.400 51.200 ;
        RECT 111.000 49.800 111.400 50.200 ;
        RECT 109.400 48.800 109.800 49.200 ;
        RECT 110.200 48.800 110.600 49.200 ;
        RECT 109.400 48.200 109.700 48.800 ;
        RECT 105.400 47.800 105.800 48.200 ;
        RECT 108.600 47.800 109.000 48.200 ;
        RECT 109.400 47.800 109.800 48.200 ;
        RECT 100.600 46.800 101.000 47.200 ;
        RECT 103.800 46.800 104.200 47.200 ;
        RECT 104.600 46.800 105.000 47.200 ;
        RECT 100.600 37.200 100.900 46.800 ;
        RECT 103.000 45.800 103.400 46.200 ;
        RECT 103.000 45.200 103.300 45.800 ;
        RECT 103.000 44.800 103.400 45.200 ;
        RECT 103.800 43.800 104.200 44.200 ;
        RECT 100.600 36.800 101.000 37.200 ;
        RECT 103.800 35.200 104.100 43.800 ;
        RECT 104.600 39.200 104.900 46.800 ;
        RECT 105.400 46.200 105.700 47.800 ;
        RECT 111.000 47.200 111.300 49.800 ;
        RECT 114.200 48.800 114.600 49.200 ;
        RECT 107.000 47.100 107.400 47.200 ;
        RECT 107.800 47.100 108.200 47.200 ;
        RECT 107.000 46.800 108.200 47.100 ;
        RECT 111.000 46.800 111.400 47.200 ;
        RECT 111.800 47.100 112.200 47.200 ;
        RECT 112.600 47.100 113.000 47.200 ;
        RECT 111.800 46.800 113.000 47.100 ;
        RECT 114.200 46.200 114.500 48.800 ;
        RECT 115.000 47.200 115.300 50.800 ;
        RECT 115.000 46.800 115.400 47.200 ;
        RECT 115.800 46.200 116.100 53.800 ;
        RECT 116.600 52.800 117.000 53.200 ;
        RECT 117.400 53.100 117.800 53.200 ;
        RECT 118.200 53.100 118.600 53.200 ;
        RECT 117.400 52.800 118.600 53.100 ;
        RECT 116.600 49.200 116.900 52.800 ;
        RECT 117.400 51.800 117.800 52.200 ;
        RECT 121.400 52.100 121.800 57.900 ;
        RECT 123.800 54.800 124.200 55.200 ;
        RECT 123.800 54.200 124.100 54.800 ;
        RECT 124.600 54.200 124.900 64.800 ;
        RECT 127.000 63.100 127.400 68.900 ;
        RECT 129.400 68.200 129.700 71.800 ;
        RECT 127.800 66.800 128.200 67.200 ;
        RECT 127.800 62.200 128.100 66.800 ;
        RECT 128.600 65.100 129.000 67.900 ;
        RECT 129.400 67.800 129.800 68.200 ;
        RECT 129.400 66.800 129.800 67.200 ;
        RECT 130.200 67.100 130.500 74.800 ;
        RECT 131.000 73.200 131.300 76.800 ;
        RECT 135.000 76.200 135.300 88.800 ;
        RECT 136.600 87.800 137.000 88.200 ;
        RECT 135.800 81.800 136.200 82.200 ;
        RECT 135.800 76.200 136.100 81.800 ;
        RECT 132.600 75.800 133.000 76.200 ;
        RECT 135.000 75.800 135.400 76.200 ;
        RECT 135.800 75.800 136.200 76.200 ;
        RECT 132.600 75.200 132.900 75.800 ;
        RECT 132.600 74.800 133.000 75.200 ;
        RECT 135.000 74.200 135.300 75.800 ;
        RECT 135.800 74.800 136.200 75.200 ;
        RECT 135.000 73.800 135.400 74.200 ;
        RECT 131.000 72.800 131.400 73.200 ;
        RECT 134.200 73.100 134.600 73.200 ;
        RECT 135.000 73.100 135.400 73.200 ;
        RECT 134.200 72.800 135.400 73.100 ;
        RECT 132.600 67.800 133.000 68.200 ;
        RECT 134.200 68.100 134.600 68.200 ;
        RECT 135.000 68.100 135.400 68.200 ;
        RECT 134.200 67.800 135.400 68.100 ;
        RECT 132.600 67.200 132.900 67.800 ;
        RECT 131.000 67.100 131.400 67.200 ;
        RECT 130.200 66.800 131.400 67.100 ;
        RECT 132.600 66.800 133.000 67.200 ;
        RECT 127.800 61.800 128.200 62.200 ;
        RECT 123.800 53.800 124.200 54.200 ;
        RECT 124.600 53.800 125.000 54.200 ;
        RECT 117.400 51.200 117.700 51.800 ;
        RECT 117.400 50.800 117.800 51.200 ;
        RECT 122.200 50.800 122.600 51.200 ;
        RECT 117.400 49.800 117.800 50.200 ;
        RECT 116.600 48.800 117.000 49.200 ;
        RECT 117.400 48.200 117.700 49.800 ;
        RECT 117.400 47.800 117.800 48.200 ;
        RECT 105.400 45.800 105.800 46.200 ;
        RECT 106.200 46.100 106.600 46.200 ;
        RECT 107.000 46.100 107.400 46.200 ;
        RECT 106.200 45.800 107.400 46.100 ;
        RECT 111.800 46.100 112.200 46.200 ;
        RECT 112.600 46.100 113.000 46.200 ;
        RECT 111.800 45.800 113.000 46.100 ;
        RECT 114.200 45.800 114.600 46.200 ;
        RECT 115.800 45.800 116.200 46.200 ;
        RECT 105.400 43.200 105.700 45.800 ;
        RECT 105.400 42.800 105.800 43.200 ;
        RECT 104.600 38.800 105.000 39.200 ;
        RECT 103.800 34.800 104.200 35.200 ;
        RECT 105.400 34.800 105.800 35.200 ;
        RECT 105.400 34.200 105.700 34.800 ;
        RECT 99.800 33.800 100.200 34.200 ;
        RECT 105.400 33.800 105.800 34.200 ;
        RECT 106.200 33.800 106.600 34.200 ;
        RECT 99.000 32.800 99.400 33.200 ;
        RECT 100.600 32.800 101.000 33.200 ;
        RECT 100.600 32.200 100.900 32.800 ;
        RECT 106.200 32.200 106.500 33.800 ;
        RECT 99.000 31.800 99.400 32.200 ;
        RECT 100.600 31.800 101.000 32.200 ;
        RECT 103.800 31.800 104.200 32.200 ;
        RECT 105.400 31.800 105.800 32.200 ;
        RECT 106.200 31.800 106.600 32.200 ;
        RECT 86.200 29.100 86.600 29.200 ;
        RECT 86.200 28.800 88.100 29.100 ;
        RECT 87.800 28.200 88.100 28.800 ;
        RECT 85.400 27.800 85.800 28.200 ;
        RECT 87.000 27.800 87.400 28.200 ;
        RECT 87.800 27.800 88.200 28.200 ;
        RECT 95.000 27.800 95.400 28.200 ;
        RECT 83.000 26.800 83.400 27.200 ;
        RECT 83.800 26.800 84.200 27.200 ;
        RECT 84.600 26.800 85.000 27.200 ;
        RECT 86.200 26.800 86.600 27.200 ;
        RECT 81.400 25.800 81.800 26.200 ;
        RECT 82.200 25.800 82.600 26.200 ;
        RECT 83.000 25.800 83.400 26.200 ;
        RECT 81.400 23.200 81.700 25.800 ;
        RECT 81.400 22.800 81.800 23.200 ;
        RECT 81.400 19.800 81.800 20.200 ;
        RECT 81.400 15.200 81.700 19.800 ;
        RECT 83.000 19.200 83.300 25.800 ;
        RECT 86.200 25.200 86.500 26.800 ;
        RECT 87.000 26.200 87.300 27.800 ;
        RECT 95.000 27.200 95.300 27.800 ;
        RECT 91.000 27.100 91.400 27.200 ;
        RECT 91.800 27.100 92.200 27.200 ;
        RECT 91.000 26.800 92.200 27.100 ;
        RECT 93.400 27.100 93.800 27.200 ;
        RECT 94.200 27.100 94.600 27.200 ;
        RECT 93.400 26.800 94.600 27.100 ;
        RECT 95.000 26.800 95.400 27.200 ;
        RECT 96.600 26.800 97.000 27.200 ;
        RECT 97.400 26.800 97.800 27.200 ;
        RECT 98.200 26.800 98.600 27.200 ;
        RECT 87.000 25.800 87.400 26.200 ;
        RECT 87.800 25.800 88.200 26.200 ;
        RECT 88.600 25.800 89.000 26.200 ;
        RECT 89.400 26.100 89.800 26.200 ;
        RECT 90.200 26.100 90.600 26.200 ;
        RECT 89.400 25.800 90.600 26.100 ;
        RECT 92.600 26.100 93.000 26.200 ;
        RECT 93.400 26.100 93.800 26.200 ;
        RECT 92.600 25.800 93.800 26.100 ;
        RECT 95.800 25.800 96.200 26.200 ;
        RECT 87.800 25.200 88.100 25.800 ;
        RECT 86.200 24.800 86.600 25.200 ;
        RECT 87.800 24.800 88.200 25.200 ;
        RECT 87.000 21.800 87.400 22.200 ;
        RECT 83.000 18.800 83.400 19.200 ;
        RECT 85.400 16.100 85.800 16.200 ;
        RECT 86.200 16.100 86.600 16.200 ;
        RECT 85.400 15.800 86.600 16.100 ;
        RECT 81.400 14.800 81.800 15.200 ;
        RECT 81.400 14.100 81.800 14.200 ;
        RECT 82.200 14.100 82.600 14.200 ;
        RECT 81.400 13.800 82.600 14.100 ;
        RECT 83.800 13.800 84.200 14.200 ;
        RECT 82.200 12.800 82.600 13.200 ;
        RECT 78.200 7.800 78.600 8.200 ;
        RECT 80.600 7.800 81.000 8.200 ;
        RECT 80.600 7.200 80.900 7.800 ;
        RECT 82.200 7.200 82.500 12.800 ;
        RECT 83.800 10.200 84.100 13.800 ;
        RECT 86.200 11.800 86.600 12.200 ;
        RECT 83.800 9.800 84.200 10.200 ;
        RECT 80.600 6.800 81.000 7.200 ;
        RECT 82.200 6.800 82.600 7.200 ;
        RECT 78.200 5.100 78.600 5.200 ;
        RECT 79.000 5.100 79.400 5.200 ;
        RECT 78.200 4.800 79.400 5.100 ;
        RECT 83.800 3.100 84.200 8.900 ;
        RECT 84.600 6.800 85.000 7.200 ;
        RECT 84.600 6.200 84.900 6.800 ;
        RECT 86.200 6.200 86.500 11.800 ;
        RECT 87.000 6.200 87.300 21.800 ;
        RECT 87.800 15.800 88.200 16.200 ;
        RECT 87.800 15.200 88.100 15.800 ;
        RECT 87.800 14.800 88.200 15.200 ;
        RECT 88.600 14.200 88.900 25.800 ;
        RECT 90.200 25.200 90.500 25.800 ;
        RECT 90.200 24.800 90.600 25.200 ;
        RECT 94.200 24.800 94.600 25.200 ;
        RECT 94.200 22.200 94.500 24.800 ;
        RECT 89.400 21.800 89.800 22.200 ;
        RECT 94.200 21.800 94.600 22.200 ;
        RECT 89.400 21.200 89.700 21.800 ;
        RECT 89.400 20.800 89.800 21.200 ;
        RECT 94.200 20.800 94.600 21.200 ;
        RECT 88.600 14.100 89.000 14.200 ;
        RECT 87.800 13.800 89.000 14.100 ;
        RECT 87.800 9.200 88.100 13.800 ;
        RECT 89.400 13.100 89.800 15.900 ;
        RECT 91.000 12.100 91.400 17.900 ;
        RECT 94.200 15.200 94.500 20.800 ;
        RECT 95.800 19.200 96.100 25.800 ;
        RECT 96.600 25.100 96.900 26.800 ;
        RECT 97.400 26.200 97.700 26.800 ;
        RECT 98.200 26.200 98.500 26.800 ;
        RECT 99.000 26.200 99.300 31.800 ;
        RECT 97.400 25.800 97.800 26.200 ;
        RECT 98.200 25.800 98.600 26.200 ;
        RECT 99.000 25.800 99.400 26.200 ;
        RECT 100.600 26.100 101.000 26.200 ;
        RECT 101.400 26.100 101.800 26.200 ;
        RECT 100.600 25.800 101.800 26.100 ;
        RECT 97.400 25.100 97.800 25.200 ;
        RECT 96.600 24.800 97.800 25.100 ;
        RECT 99.000 19.200 99.300 25.800 ;
        RECT 100.600 21.800 101.000 22.200 ;
        RECT 100.600 21.200 100.900 21.800 ;
        RECT 100.600 20.800 101.000 21.200 ;
        RECT 95.800 18.800 96.200 19.200 ;
        RECT 99.000 18.800 99.400 19.200 ;
        RECT 94.200 14.800 94.600 15.200 ;
        RECT 91.800 12.800 92.200 13.200 ;
        RECT 91.000 9.800 91.400 10.200 ;
        RECT 91.000 9.200 91.300 9.800 ;
        RECT 87.800 8.800 88.200 9.200 ;
        RECT 84.600 5.800 85.000 6.200 ;
        RECT 86.200 5.800 86.600 6.200 ;
        RECT 87.000 5.800 87.400 6.200 ;
        RECT 88.600 3.100 89.000 8.900 ;
        RECT 91.000 8.800 91.400 9.200 ;
        RECT 90.200 5.100 90.600 7.900 ;
        RECT 91.800 7.200 92.100 12.800 ;
        RECT 95.800 12.100 96.200 17.900 ;
        RECT 102.200 17.800 102.600 18.200 ;
        RECT 100.600 16.800 101.000 17.200 ;
        RECT 99.800 14.800 100.200 15.200 ;
        RECT 99.800 14.200 100.100 14.800 ;
        RECT 98.200 13.800 98.600 14.200 ;
        RECT 99.800 13.800 100.200 14.200 ;
        RECT 98.200 13.200 98.500 13.800 ;
        RECT 100.600 13.200 100.900 16.800 ;
        RECT 102.200 15.200 102.500 17.800 ;
        RECT 102.200 14.800 102.600 15.200 ;
        RECT 98.200 12.800 98.600 13.200 ;
        RECT 99.000 13.100 99.400 13.200 ;
        RECT 99.800 13.100 100.200 13.200 ;
        RECT 99.000 12.800 100.200 13.100 ;
        RECT 100.600 12.800 101.000 13.200 ;
        RECT 103.800 9.200 104.100 31.800 ;
        RECT 105.400 29.200 105.700 31.800 ;
        RECT 105.400 28.800 105.800 29.200 ;
        RECT 104.600 27.800 105.000 28.200 ;
        RECT 104.600 27.200 104.900 27.800 ;
        RECT 104.600 26.800 105.000 27.200 ;
        RECT 106.200 26.800 106.600 27.200 ;
        RECT 106.200 23.200 106.500 26.800 ;
        RECT 107.000 26.200 107.300 45.800 ;
        RECT 112.600 45.100 113.000 45.200 ;
        RECT 113.400 45.100 113.800 45.200 ;
        RECT 112.600 44.800 113.800 45.100 ;
        RECT 114.200 44.800 114.600 45.200 ;
        RECT 111.000 39.800 111.400 40.200 ;
        RECT 108.600 37.100 109.000 37.200 ;
        RECT 109.400 37.100 109.800 37.200 ;
        RECT 108.600 36.800 109.800 37.100 ;
        RECT 111.000 35.200 111.300 39.800 ;
        RECT 111.800 36.800 112.200 37.200 ;
        RECT 111.800 35.200 112.100 36.800 ;
        RECT 107.800 34.800 108.200 35.200 ;
        RECT 110.200 34.800 110.600 35.200 ;
        RECT 111.000 34.800 111.400 35.200 ;
        RECT 111.800 34.800 112.200 35.200 ;
        RECT 107.800 29.200 108.100 34.800 ;
        RECT 110.200 34.200 110.500 34.800 ;
        RECT 110.200 33.800 110.600 34.200 ;
        RECT 111.800 31.200 112.100 34.800 ;
        RECT 112.600 34.100 113.000 34.200 ;
        RECT 113.400 34.100 113.800 34.200 ;
        RECT 112.600 33.800 113.800 34.100 ;
        RECT 114.200 33.200 114.500 44.800 ;
        RECT 120.600 43.100 121.000 48.900 ;
        RECT 122.200 46.200 122.500 50.800 ;
        RECT 124.600 48.200 124.900 53.800 ;
        RECT 126.200 52.100 126.600 57.900 ;
        RECT 127.800 53.100 128.200 55.900 ;
        RECT 129.400 55.200 129.700 66.800 ;
        RECT 135.800 66.200 136.100 74.800 ;
        RECT 136.600 74.200 136.900 87.800 ;
        RECT 139.800 83.100 140.200 88.900 ;
        RECT 142.200 88.200 142.500 94.800 ;
        RECT 144.600 94.200 144.900 98.800 ;
        RECT 147.000 95.800 147.400 96.200 ;
        RECT 145.400 94.800 145.800 95.200 ;
        RECT 145.400 94.200 145.700 94.800 ;
        RECT 147.000 94.200 147.300 95.800 ;
        RECT 147.800 94.800 148.200 95.200 ;
        RECT 143.800 93.800 144.200 94.200 ;
        RECT 144.600 93.800 145.000 94.200 ;
        RECT 145.400 93.800 145.800 94.200 ;
        RECT 147.000 93.800 147.400 94.200 ;
        RECT 143.800 93.200 144.100 93.800 ;
        RECT 147.800 93.200 148.100 94.800 ;
        RECT 148.600 94.200 148.900 98.800 ;
        RECT 151.800 98.200 152.100 112.800 ;
        RECT 152.600 103.100 153.000 108.900 ;
        RECT 154.200 103.200 154.500 112.800 ;
        RECT 155.800 112.200 156.100 112.800 ;
        RECT 158.200 112.200 158.500 112.800 ;
        RECT 159.000 112.200 159.300 112.800 ;
        RECT 155.800 111.800 156.200 112.200 ;
        RECT 158.200 111.800 158.600 112.200 ;
        RECT 159.000 111.800 159.400 112.200 ;
        RECT 163.800 111.800 164.200 112.200 ;
        RECT 155.800 109.800 156.200 110.200 ;
        RECT 162.200 109.800 162.600 110.200 ;
        RECT 155.800 106.200 156.100 109.800 ;
        RECT 162.200 109.200 162.500 109.800 ;
        RECT 155.800 105.800 156.200 106.200 ;
        RECT 154.200 102.800 154.600 103.200 ;
        RECT 157.400 103.100 157.800 108.900 ;
        RECT 159.800 108.800 160.200 109.200 ;
        RECT 162.200 108.800 162.600 109.200 ;
        RECT 159.800 108.200 160.100 108.800 ;
        RECT 159.800 107.800 160.200 108.200 ;
        RECT 163.800 107.200 164.100 111.800 ;
        RECT 164.600 108.100 165.000 108.200 ;
        RECT 165.400 108.100 165.800 108.200 ;
        RECT 164.600 107.800 165.800 108.100 ;
        RECT 160.600 107.100 161.000 107.200 ;
        RECT 161.400 107.100 161.800 107.200 ;
        RECT 160.600 106.800 161.800 107.100 ;
        RECT 163.800 106.800 164.200 107.200 ;
        RECT 163.800 106.200 164.100 106.800 ;
        RECT 166.200 106.200 166.500 115.800 ;
        RECT 160.600 105.800 161.000 106.200 ;
        RECT 163.800 105.800 164.200 106.200 ;
        RECT 165.400 106.100 165.800 106.200 ;
        RECT 166.200 106.100 166.600 106.200 ;
        RECT 165.400 105.800 166.600 106.100 ;
        RECT 160.600 103.200 160.900 105.800 ;
        RECT 160.600 102.800 161.000 103.200 ;
        RECT 151.800 97.800 152.200 98.200 ;
        RECT 151.000 94.800 151.400 95.200 ;
        RECT 151.000 94.200 151.300 94.800 ;
        RECT 148.600 93.800 149.000 94.200 ;
        RECT 149.400 94.100 149.800 94.200 ;
        RECT 150.200 94.100 150.600 94.200 ;
        RECT 149.400 93.800 150.600 94.100 ;
        RECT 151.000 93.800 151.400 94.200 ;
        RECT 151.800 94.100 152.100 97.800 ;
        RECT 161.400 96.800 161.800 97.200 ;
        RECT 161.400 95.200 161.700 96.800 ;
        RECT 163.000 96.100 163.400 96.200 ;
        RECT 163.800 96.100 164.200 96.200 ;
        RECT 163.000 95.800 164.200 96.100 ;
        RECT 166.200 95.800 166.600 96.200 ;
        RECT 156.600 94.800 157.000 95.200 ;
        RECT 161.400 94.800 161.800 95.200 ;
        RECT 152.600 94.100 153.000 94.200 ;
        RECT 151.800 93.800 153.000 94.100 ;
        RECT 143.800 92.800 144.200 93.200 ;
        RECT 147.800 92.800 148.200 93.200 ;
        RECT 147.000 91.800 147.400 92.200 ;
        RECT 147.000 90.200 147.300 91.800 ;
        RECT 147.000 89.800 147.400 90.200 ;
        RECT 142.200 87.800 142.600 88.200 ;
        RECT 143.800 86.800 144.200 87.200 ;
        RECT 143.800 86.300 144.100 86.800 ;
        RECT 143.800 85.900 144.200 86.300 ;
        RECT 144.600 83.100 145.000 88.900 ;
        RECT 145.400 86.800 145.800 87.200 ;
        RECT 145.400 86.200 145.700 86.800 ;
        RECT 145.400 85.800 145.800 86.200 ;
        RECT 146.200 85.100 146.600 87.900 ;
        RECT 148.600 87.100 148.900 93.800 ;
        RECT 152.600 93.200 152.900 93.800 ;
        RECT 150.200 93.100 150.600 93.200 ;
        RECT 151.000 93.100 151.400 93.200 ;
        RECT 150.200 92.800 151.400 93.100 ;
        RECT 152.600 92.800 153.000 93.200 ;
        RECT 154.200 93.100 154.600 93.200 ;
        RECT 155.000 93.100 155.400 93.200 ;
        RECT 154.200 92.800 155.400 93.100 ;
        RECT 150.200 90.800 150.600 91.200 ;
        RECT 150.200 89.200 150.500 90.800 ;
        RECT 150.200 88.800 150.600 89.200 ;
        RECT 151.800 88.800 152.200 89.200 ;
        RECT 149.400 87.100 149.800 87.200 ;
        RECT 148.600 86.800 149.800 87.100 ;
        RECT 150.200 86.200 150.500 88.800 ;
        RECT 151.800 86.200 152.100 88.800 ;
        RECT 156.600 88.200 156.900 94.800 ;
        RECT 157.400 93.800 157.800 94.200 ;
        RECT 160.600 93.800 161.000 94.200 ;
        RECT 161.400 93.800 161.800 94.200 ;
        RECT 157.400 89.200 157.700 93.800 ;
        RECT 160.600 93.200 160.900 93.800 ;
        RECT 159.000 93.100 159.400 93.200 ;
        RECT 159.800 93.100 160.200 93.200 ;
        RECT 159.000 92.800 160.200 93.100 ;
        RECT 160.600 92.800 161.000 93.200 ;
        RECT 161.400 92.200 161.700 93.800 ;
        RECT 161.400 91.800 161.800 92.200 ;
        RECT 163.800 90.200 164.100 95.800 ;
        RECT 166.200 95.200 166.500 95.800 ;
        RECT 167.000 95.200 167.300 115.800 ;
        RECT 169.400 115.200 169.700 116.800 ;
        RECT 169.400 114.800 169.800 115.200 ;
        RECT 171.800 112.100 172.200 118.900 ;
        RECT 172.600 112.100 173.000 118.900 ;
        RECT 173.400 112.100 173.800 117.900 ;
        RECT 174.200 114.200 174.500 123.800 ;
        RECT 175.800 121.800 176.200 122.200 ;
        RECT 180.600 121.800 181.000 122.200 ;
        RECT 188.600 121.800 189.000 122.200 ;
        RECT 191.000 121.800 191.400 122.200 ;
        RECT 174.200 113.800 174.600 114.200 ;
        RECT 175.000 112.100 175.400 117.900 ;
        RECT 175.800 116.200 176.100 121.800 ;
        RECT 175.800 115.800 176.200 116.200 ;
        RECT 175.800 113.800 176.200 114.200 ;
        RECT 175.800 113.200 176.100 113.800 ;
        RECT 175.800 112.800 176.200 113.200 ;
        RECT 176.600 112.100 177.000 117.900 ;
        RECT 177.400 112.100 177.800 118.900 ;
        RECT 178.200 112.100 178.600 118.900 ;
        RECT 179.000 112.100 179.400 118.900 ;
        RECT 167.800 108.800 168.200 109.200 ;
        RECT 171.000 108.800 171.400 109.200 ;
        RECT 172.600 109.100 173.000 109.200 ;
        RECT 173.400 109.100 173.800 109.200 ;
        RECT 172.600 108.800 173.800 109.100 ;
        RECT 167.800 108.200 168.100 108.800 ;
        RECT 171.000 108.200 171.300 108.800 ;
        RECT 167.800 107.800 168.200 108.200 ;
        RECT 168.600 108.100 169.000 108.200 ;
        RECT 169.400 108.100 169.800 108.200 ;
        RECT 168.600 107.800 169.800 108.100 ;
        RECT 171.000 107.800 171.400 108.200 ;
        RECT 175.000 107.800 175.400 108.200 ;
        RECT 175.800 108.100 176.200 108.200 ;
        RECT 176.600 108.100 177.000 108.200 ;
        RECT 175.800 107.800 177.000 108.100 ;
        RECT 171.000 106.200 171.300 107.800 ;
        RECT 175.000 107.200 175.300 107.800 ;
        RECT 175.000 106.800 175.400 107.200 ;
        RECT 169.400 105.800 169.800 106.200 ;
        RECT 170.200 105.800 170.600 106.200 ;
        RECT 171.000 105.800 171.400 106.200 ;
        RECT 172.600 105.800 173.000 106.200 ;
        RECT 169.400 100.200 169.700 105.800 ;
        RECT 169.400 99.800 169.800 100.200 ;
        RECT 167.800 97.800 168.200 98.200 ;
        RECT 167.800 96.200 168.100 97.800 ;
        RECT 167.800 95.800 168.200 96.200 ;
        RECT 169.400 95.800 169.800 96.200 ;
        RECT 166.200 94.800 166.600 95.200 ;
        RECT 167.000 94.800 167.400 95.200 ;
        RECT 166.200 94.100 166.600 94.200 ;
        RECT 167.000 94.100 167.400 94.200 ;
        RECT 166.200 93.800 167.400 94.100 ;
        RECT 167.800 93.200 168.100 95.800 ;
        RECT 169.400 95.200 169.700 95.800 ;
        RECT 169.400 94.800 169.800 95.200 ;
        RECT 170.200 94.200 170.500 105.800 ;
        RECT 172.600 105.200 172.900 105.800 ;
        RECT 172.600 105.100 173.000 105.200 ;
        RECT 172.600 104.800 173.700 105.100 ;
        RECT 171.800 96.800 172.200 97.200 ;
        RECT 171.800 96.200 172.100 96.800 ;
        RECT 171.800 95.800 172.200 96.200 ;
        RECT 171.800 95.100 172.200 95.200 ;
        RECT 171.800 94.800 172.900 95.100 ;
        RECT 170.200 93.800 170.600 94.200 ;
        RECT 171.000 93.800 171.400 94.200 ;
        RECT 167.800 92.800 168.200 93.200 ;
        RECT 164.600 91.800 165.000 92.200 ;
        RECT 167.800 91.800 168.200 92.200 ;
        RECT 158.200 89.800 158.600 90.200 ;
        RECT 163.800 89.800 164.200 90.200 ;
        RECT 157.400 88.800 157.800 89.200 ;
        RECT 156.600 88.100 157.000 88.200 ;
        RECT 155.800 87.800 157.000 88.100 ;
        RECT 148.600 86.100 149.000 86.200 ;
        RECT 149.400 86.100 149.800 86.200 ;
        RECT 148.600 85.800 149.800 86.100 ;
        RECT 150.200 85.800 150.600 86.200 ;
        RECT 151.000 86.100 151.400 86.200 ;
        RECT 151.800 86.100 152.200 86.200 ;
        RECT 151.000 85.800 152.200 86.100 ;
        RECT 153.400 85.800 153.800 86.200 ;
        RECT 147.000 85.100 147.400 85.200 ;
        RECT 147.800 85.100 148.200 85.200 ;
        RECT 147.000 84.800 148.200 85.100 ;
        RECT 147.000 83.800 147.400 84.200 ;
        RECT 137.400 76.800 137.800 77.200 ;
        RECT 139.800 76.800 140.200 77.200 ;
        RECT 141.400 76.800 141.800 77.200 ;
        RECT 137.400 75.200 137.700 76.800 ;
        RECT 139.800 76.200 140.100 76.800 ;
        RECT 139.800 75.800 140.200 76.200 ;
        RECT 137.400 74.800 137.800 75.200 ;
        RECT 141.400 74.200 141.700 76.800 ;
        RECT 136.600 73.800 137.000 74.200 ;
        RECT 141.400 73.800 141.800 74.200 ;
        RECT 136.600 72.200 136.900 73.800 ;
        RECT 139.000 73.100 139.400 73.200 ;
        RECT 139.800 73.100 140.200 73.200 ;
        RECT 142.200 73.100 142.600 75.900 ;
        RECT 143.000 73.800 143.400 74.200 ;
        RECT 143.000 73.200 143.300 73.800 ;
        RECT 139.000 72.800 140.200 73.100 ;
        RECT 143.000 72.800 143.400 73.200 ;
        RECT 136.600 71.800 137.000 72.200 ;
        RECT 143.800 72.100 144.200 77.900 ;
        RECT 144.600 74.700 145.000 75.100 ;
        RECT 144.600 74.200 144.900 74.700 ;
        RECT 144.600 73.800 145.000 74.200 ;
        RECT 136.600 67.200 136.900 71.800 ;
        RECT 139.800 69.800 140.200 70.200 ;
        RECT 141.400 69.800 141.800 70.200 ;
        RECT 139.800 69.200 140.100 69.800 ;
        RECT 139.800 68.800 140.200 69.200 ;
        RECT 140.600 68.800 141.000 69.200 ;
        RECT 140.600 68.200 140.900 68.800 ;
        RECT 140.600 67.800 141.000 68.200 ;
        RECT 136.600 66.800 137.000 67.200 ;
        RECT 137.400 66.800 137.800 67.200 ;
        RECT 139.000 66.800 139.400 67.200 ;
        RECT 137.400 66.200 137.700 66.800 ;
        RECT 130.200 66.100 130.600 66.200 ;
        RECT 131.000 66.100 131.400 66.200 ;
        RECT 130.200 65.800 131.400 66.100 ;
        RECT 132.600 65.800 133.000 66.200 ;
        RECT 135.800 65.800 136.200 66.200 ;
        RECT 136.600 65.800 137.000 66.200 ;
        RECT 137.400 65.800 137.800 66.200 ;
        RECT 138.200 65.800 138.600 66.200 ;
        RECT 131.800 64.800 132.200 65.200 ;
        RECT 131.800 56.200 132.100 64.800 ;
        RECT 130.200 55.800 130.600 56.200 ;
        RECT 131.800 55.800 132.200 56.200 ;
        RECT 130.200 55.200 130.500 55.800 ;
        RECT 129.400 54.800 129.800 55.200 ;
        RECT 130.200 54.800 130.600 55.200 ;
        RECT 131.800 54.200 132.100 55.800 ;
        RECT 128.600 54.100 129.000 54.200 ;
        RECT 129.400 54.100 129.800 54.200 ;
        RECT 128.600 53.800 129.800 54.100 ;
        RECT 131.800 53.800 132.200 54.200 ;
        RECT 124.600 47.800 125.000 48.200 ;
        RECT 122.200 45.800 122.600 46.200 ;
        RECT 122.200 42.800 122.600 43.200 ;
        RECT 125.400 43.100 125.800 48.900 ;
        RECT 126.200 46.800 126.600 47.200 ;
        RECT 126.200 45.200 126.500 46.800 ;
        RECT 126.200 44.800 126.600 45.200 ;
        RECT 127.000 45.100 127.400 47.900 ;
        RECT 127.800 46.800 128.200 47.200 ;
        RECT 127.800 46.200 128.100 46.800 ;
        RECT 127.800 45.800 128.200 46.200 ;
        RECT 127.800 44.800 128.200 45.200 ;
        RECT 127.800 44.200 128.100 44.800 ;
        RECT 127.800 43.800 128.200 44.200 ;
        RECT 115.000 34.100 115.400 34.200 ;
        RECT 115.800 34.100 116.200 34.200 ;
        RECT 115.000 33.800 116.200 34.100 ;
        RECT 114.200 32.800 114.600 33.200 ;
        RECT 115.800 32.800 116.200 33.200 ;
        RECT 112.600 31.800 113.000 32.200 ;
        RECT 113.400 31.800 113.800 32.200 ;
        RECT 111.800 30.800 112.200 31.200 ;
        RECT 107.800 28.800 108.200 29.200 ;
        RECT 107.000 25.800 107.400 26.200 ;
        RECT 104.600 22.800 105.000 23.200 ;
        RECT 106.200 22.800 106.600 23.200 ;
        RECT 104.600 19.200 104.900 22.800 ;
        RECT 104.600 18.800 105.000 19.200 ;
        RECT 107.000 12.100 107.400 17.900 ;
        RECT 102.200 9.100 102.600 9.200 ;
        RECT 103.000 9.100 103.400 9.200 ;
        RECT 91.800 6.800 92.200 7.200 ;
        RECT 93.400 3.100 93.800 8.900 ;
        RECT 94.200 6.800 94.600 7.200 ;
        RECT 94.200 6.200 94.500 6.800 ;
        RECT 94.200 5.800 94.600 6.200 ;
        RECT 95.800 6.100 96.200 6.200 ;
        RECT 96.600 6.100 97.000 6.200 ;
        RECT 95.800 5.800 97.000 6.100 ;
        RECT 98.200 3.100 98.600 8.900 ;
        RECT 102.200 8.800 103.400 9.100 ;
        RECT 103.800 8.800 104.200 9.200 ;
        RECT 99.800 5.100 100.200 7.900 ;
        RECT 104.600 3.100 105.000 8.900 ;
        RECT 107.800 8.200 108.100 28.800 ;
        RECT 111.800 27.800 112.200 28.200 ;
        RECT 111.800 27.200 112.100 27.800 ;
        RECT 112.600 27.200 112.900 31.800 ;
        RECT 113.400 27.200 113.700 31.800 ;
        RECT 115.800 27.200 116.100 32.800 ;
        RECT 119.000 32.100 119.400 37.900 ;
        RECT 120.600 36.800 121.000 37.200 ;
        RECT 120.600 35.200 120.900 36.800 ;
        RECT 120.600 34.800 121.000 35.200 ;
        RECT 119.000 29.800 119.400 30.200 ;
        RECT 119.000 27.200 119.300 29.800 ;
        RECT 121.400 27.800 121.800 28.200 ;
        RECT 109.400 26.800 109.800 27.200 ;
        RECT 111.800 26.800 112.200 27.200 ;
        RECT 112.600 26.800 113.000 27.200 ;
        RECT 113.400 26.800 113.800 27.200 ;
        RECT 115.800 26.800 116.200 27.200 ;
        RECT 116.600 26.800 117.000 27.200 ;
        RECT 119.000 26.800 119.400 27.200 ;
        RECT 109.400 26.200 109.700 26.800 ;
        RECT 109.400 25.800 109.800 26.200 ;
        RECT 112.600 25.800 113.000 26.200 ;
        RECT 113.400 25.800 113.800 26.200 ;
        RECT 115.000 25.800 115.400 26.200 ;
        RECT 112.600 25.200 112.900 25.800 ;
        RECT 113.400 25.200 113.700 25.800 ;
        RECT 112.600 24.800 113.000 25.200 ;
        RECT 113.400 24.800 113.800 25.200 ;
        RECT 110.200 21.800 110.600 22.200 ;
        RECT 110.200 15.200 110.500 21.800 ;
        RECT 110.200 14.800 110.600 15.200 ;
        RECT 110.200 13.800 110.600 14.200 ;
        RECT 110.200 12.200 110.500 13.800 ;
        RECT 110.200 11.800 110.600 12.200 ;
        RECT 111.800 12.100 112.200 17.900 ;
        RECT 115.000 17.200 115.300 25.800 ;
        RECT 115.800 21.200 116.100 26.800 ;
        RECT 116.600 25.200 116.900 26.800 ;
        RECT 121.400 26.200 121.700 27.800 ;
        RECT 122.200 27.200 122.500 42.800 ;
        RECT 124.600 39.800 125.000 40.200 ;
        RECT 123.800 32.100 124.200 37.900 ;
        RECT 124.600 34.200 124.900 39.800 ;
        RECT 128.600 39.200 128.900 53.800 ;
        RECT 129.400 51.800 129.800 52.200 ;
        RECT 129.400 46.200 129.700 51.800 ;
        RECT 132.600 51.200 132.900 65.800 ;
        RECT 133.400 65.100 133.800 65.200 ;
        RECT 134.200 65.100 134.600 65.200 ;
        RECT 133.400 64.800 134.600 65.100 ;
        RECT 135.000 61.800 135.400 62.200 ;
        RECT 133.400 54.800 133.800 55.200 ;
        RECT 133.400 54.200 133.700 54.800 ;
        RECT 133.400 53.800 133.800 54.200 ;
        RECT 133.400 52.800 133.800 53.200 ;
        RECT 134.200 53.100 134.600 55.900 ;
        RECT 135.000 54.200 135.300 61.800 ;
        RECT 136.600 59.200 136.900 65.800 ;
        RECT 137.400 65.200 137.700 65.800 ;
        RECT 137.400 64.800 137.800 65.200 ;
        RECT 136.600 58.800 137.000 59.200 ;
        RECT 135.000 53.800 135.400 54.200 ;
        RECT 132.600 50.800 133.000 51.200 ;
        RECT 133.400 48.200 133.700 52.800 ;
        RECT 135.800 52.100 136.200 57.900 ;
        RECT 136.600 55.800 137.000 56.200 ;
        RECT 136.600 55.100 136.900 55.800 ;
        RECT 136.600 54.700 137.000 55.100 ;
        RECT 134.200 49.100 134.600 49.200 ;
        RECT 135.000 49.100 135.400 49.200 ;
        RECT 134.200 48.800 135.400 49.100 ;
        RECT 133.400 47.800 133.800 48.200 ;
        RECT 130.200 46.800 130.600 47.200 ;
        RECT 130.200 46.200 130.500 46.800 ;
        RECT 133.400 46.200 133.700 47.800 ;
        RECT 129.400 45.800 129.800 46.200 ;
        RECT 130.200 45.800 130.600 46.200 ;
        RECT 133.400 45.800 133.800 46.200 ;
        RECT 136.600 43.100 137.000 48.900 ;
        RECT 138.200 46.200 138.500 65.800 ;
        RECT 139.000 54.200 139.300 66.800 ;
        RECT 141.400 66.200 141.700 69.800 ;
        RECT 144.600 68.100 145.000 68.200 ;
        RECT 145.400 68.100 145.800 68.200 ;
        RECT 144.600 67.800 145.800 68.100 ;
        RECT 146.200 67.800 146.600 68.200 ;
        RECT 144.600 66.800 145.000 67.200 ;
        RECT 144.600 66.200 144.900 66.800 ;
        RECT 146.200 66.200 146.500 67.800 ;
        RECT 147.000 67.200 147.300 83.800 ;
        RECT 153.400 83.200 153.700 85.800 ;
        RECT 153.400 82.800 153.800 83.200 ;
        RECT 148.600 81.800 149.000 82.200 ;
        RECT 148.600 79.200 148.900 81.800 ;
        RECT 148.600 78.800 149.000 79.200 ;
        RECT 153.400 78.800 153.800 79.200 ;
        RECT 147.800 75.800 148.200 76.200 ;
        RECT 147.800 68.200 148.100 75.800 ;
        RECT 148.600 72.100 149.000 77.900 ;
        RECT 150.200 77.100 150.600 77.200 ;
        RECT 151.000 77.100 151.400 77.200 ;
        RECT 150.200 76.800 151.400 77.100 ;
        RECT 149.400 75.800 149.800 76.200 ;
        RECT 149.400 69.200 149.700 75.800 ;
        RECT 153.400 75.200 153.700 78.800 ;
        RECT 153.400 74.800 153.800 75.200 ;
        RECT 154.200 74.100 154.600 74.200 ;
        RECT 155.000 74.100 155.400 74.200 ;
        RECT 154.200 73.800 155.400 74.100 ;
        RECT 155.800 73.200 156.100 87.800 ;
        RECT 158.200 87.200 158.500 89.800 ;
        RECT 164.600 89.200 164.900 91.800 ;
        RECT 159.000 88.800 159.400 89.200 ;
        RECT 159.000 87.200 159.300 88.800 ;
        RECT 156.600 86.800 157.000 87.200 ;
        RECT 158.200 86.800 158.600 87.200 ;
        RECT 159.000 86.800 159.400 87.200 ;
        RECT 156.600 86.200 156.900 86.800 ;
        RECT 156.600 85.800 157.000 86.200 ;
        RECT 159.000 85.800 159.400 86.200 ;
        RECT 159.000 85.200 159.300 85.800 ;
        RECT 159.000 84.800 159.400 85.200 ;
        RECT 163.800 83.100 164.200 88.900 ;
        RECT 164.600 88.800 165.000 89.200 ;
        RECT 165.400 87.800 165.800 88.200 ;
        RECT 164.600 86.800 165.000 87.200 ;
        RECT 164.600 86.200 164.900 86.800 ;
        RECT 164.600 85.800 165.000 86.200 ;
        RECT 163.000 80.800 163.400 81.200 ;
        RECT 156.600 76.800 157.000 77.200 ;
        RECT 156.600 73.200 156.900 76.800 ;
        RECT 157.400 76.100 157.800 76.200 ;
        RECT 158.200 76.100 158.600 76.200 ;
        RECT 157.400 75.800 158.600 76.100 ;
        RECT 159.000 75.800 159.400 76.200 ;
        RECT 160.600 76.100 161.000 76.200 ;
        RECT 161.400 76.100 161.800 76.200 ;
        RECT 160.600 75.800 161.800 76.100 ;
        RECT 159.000 75.200 159.300 75.800 ;
        RECT 159.000 74.800 159.400 75.200 ;
        RECT 159.800 74.800 160.200 75.200 ;
        RECT 159.800 74.200 160.100 74.800 ;
        RECT 163.000 74.200 163.300 80.800 ;
        RECT 157.400 74.100 157.800 74.200 ;
        RECT 158.200 74.100 158.600 74.200 ;
        RECT 157.400 73.800 158.600 74.100 ;
        RECT 159.800 73.800 160.200 74.200 ;
        RECT 160.600 73.800 161.000 74.200 ;
        RECT 163.000 73.800 163.400 74.200 ;
        RECT 154.200 73.100 154.600 73.200 ;
        RECT 155.000 73.100 155.400 73.200 ;
        RECT 154.200 72.800 155.400 73.100 ;
        RECT 155.800 72.800 156.200 73.200 ;
        RECT 156.600 72.800 157.000 73.200 ;
        RECT 149.400 68.800 149.800 69.200 ;
        RECT 154.200 68.800 154.600 69.200 ;
        RECT 147.800 67.800 148.200 68.200 ;
        RECT 150.200 67.800 150.600 68.200 ;
        RECT 153.400 67.800 153.800 68.200 ;
        RECT 147.800 67.200 148.100 67.800 ;
        RECT 150.200 67.200 150.500 67.800 ;
        RECT 153.400 67.200 153.700 67.800 ;
        RECT 147.000 66.800 147.400 67.200 ;
        RECT 147.800 66.800 148.200 67.200 ;
        RECT 150.200 66.800 150.600 67.200 ;
        RECT 151.000 66.800 151.400 67.200 ;
        RECT 151.800 66.800 152.200 67.200 ;
        RECT 153.400 66.800 153.800 67.200 ;
        RECT 151.000 66.200 151.300 66.800 ;
        RECT 151.800 66.200 152.100 66.800 ;
        RECT 141.400 65.800 141.800 66.200 ;
        RECT 144.600 65.800 145.000 66.200 ;
        RECT 146.200 65.800 146.600 66.200 ;
        RECT 147.800 65.800 148.200 66.200 ;
        RECT 151.000 65.800 151.400 66.200 ;
        RECT 151.800 65.800 152.200 66.200 ;
        RECT 141.400 60.200 141.700 65.800 ;
        RECT 147.800 65.200 148.100 65.800 ;
        RECT 154.200 65.200 154.500 68.800 ;
        RECT 147.800 65.100 148.200 65.200 ;
        RECT 147.000 64.800 148.200 65.100 ;
        RECT 154.200 64.800 154.600 65.200 ;
        RECT 155.800 65.100 156.200 67.900 ;
        RECT 156.600 66.800 157.000 67.200 ;
        RECT 141.400 59.800 141.800 60.200 ;
        RECT 147.000 59.200 147.300 64.800 ;
        RECT 147.000 58.800 147.400 59.200 ;
        RECT 153.400 58.800 153.800 59.200 ;
        RECT 139.800 54.800 140.200 55.200 ;
        RECT 139.000 53.800 139.400 54.200 ;
        RECT 139.800 47.200 140.100 54.800 ;
        RECT 140.600 52.100 141.000 57.900 ;
        RECT 143.800 54.800 144.200 55.200 ;
        RECT 141.400 54.100 141.800 54.200 ;
        RECT 142.200 54.100 142.600 54.200 ;
        RECT 141.400 53.800 142.600 54.100 ;
        RECT 143.800 53.200 144.100 54.800 ;
        RECT 143.800 52.800 144.200 53.200 ;
        RECT 145.400 51.800 145.800 52.200 ;
        RECT 149.400 52.100 149.800 57.900 ;
        RECT 150.200 55.100 150.600 55.200 ;
        RECT 151.000 55.100 151.400 55.200 ;
        RECT 150.200 54.800 151.400 55.100 ;
        RECT 153.400 55.100 153.700 58.800 ;
        RECT 153.400 54.700 153.800 55.100 ;
        RECT 154.200 52.100 154.600 57.900 ;
        RECT 155.800 53.100 156.200 55.900 ;
        RECT 156.600 54.200 156.900 66.800 ;
        RECT 157.400 63.100 157.800 68.900 ;
        RECT 160.600 68.200 160.900 73.800 ;
        RECT 161.400 71.800 161.800 72.200 ;
        RECT 161.400 69.200 161.700 71.800 ;
        RECT 161.400 68.800 161.800 69.200 ;
        RECT 160.600 67.800 161.000 68.200 ;
        RECT 158.200 66.800 158.600 67.200 ;
        RECT 158.200 66.300 158.500 66.800 ;
        RECT 158.200 65.900 158.600 66.300 ;
        RECT 158.200 65.800 158.500 65.900 ;
        RECT 159.000 55.800 159.400 56.200 ;
        RECT 159.000 55.200 159.300 55.800 ;
        RECT 159.000 54.800 159.400 55.200 ;
        RECT 156.600 53.800 157.000 54.200 ;
        RECT 159.000 52.200 159.300 54.800 ;
        RECT 159.000 51.800 159.400 52.200 ;
        RECT 145.400 49.200 145.700 51.800 ;
        RECT 159.800 50.800 160.200 51.200 ;
        RECT 139.800 46.800 140.200 47.200 ;
        RECT 140.600 46.800 141.000 47.200 ;
        RECT 138.200 45.800 138.600 46.200 ;
        RECT 131.800 41.800 132.200 42.200 ;
        RECT 128.600 38.800 129.000 39.200 ;
        RECT 124.600 33.800 125.000 34.200 ;
        RECT 125.400 33.100 125.800 35.900 ;
        RECT 127.800 35.100 128.200 35.200 ;
        RECT 128.600 35.100 129.000 35.200 ;
        RECT 127.800 34.800 129.000 35.100 ;
        RECT 130.200 34.800 130.600 35.200 ;
        RECT 130.200 34.200 130.500 34.800 ;
        RECT 127.800 33.800 128.200 34.200 ;
        RECT 130.200 33.800 130.600 34.200 ;
        RECT 126.200 32.800 126.600 33.200 ;
        RECT 122.200 26.800 122.600 27.200 ;
        RECT 124.600 27.100 125.000 27.200 ;
        RECT 125.400 27.100 125.800 27.200 ;
        RECT 124.600 26.800 125.800 27.100 ;
        RECT 126.200 27.100 126.500 32.800 ;
        RECT 127.800 29.200 128.100 33.800 ;
        RECT 129.400 32.100 129.800 32.200 ;
        RECT 130.200 32.100 130.600 32.200 ;
        RECT 129.400 31.800 130.600 32.100 ;
        RECT 127.800 28.800 128.200 29.200 ;
        RECT 131.800 27.200 132.100 41.800 ;
        RECT 139.800 40.200 140.100 46.800 ;
        RECT 140.600 46.300 140.900 46.800 ;
        RECT 140.600 45.900 141.000 46.300 ;
        RECT 141.400 43.100 141.800 48.900 ;
        RECT 143.800 48.800 144.200 49.200 ;
        RECT 145.400 48.800 145.800 49.200 ;
        RECT 151.800 48.800 152.200 49.200 ;
        RECT 143.800 48.200 144.100 48.800 ;
        RECT 143.000 45.100 143.400 47.900 ;
        RECT 143.800 47.800 144.200 48.200 ;
        RECT 147.800 47.800 148.200 48.200 ;
        RECT 149.400 48.100 149.800 48.200 ;
        RECT 150.200 48.100 150.600 48.200 ;
        RECT 149.400 47.800 150.600 48.100 ;
        RECT 147.800 47.200 148.100 47.800 ;
        RECT 151.800 47.200 152.100 48.800 ;
        RECT 159.800 47.200 160.100 50.800 ;
        RECT 145.400 46.800 145.800 47.200 ;
        RECT 146.200 46.800 146.600 47.200 ;
        RECT 147.800 46.800 148.200 47.200 ;
        RECT 148.600 46.800 149.000 47.200 ;
        RECT 151.800 46.800 152.200 47.200 ;
        RECT 159.800 46.800 160.200 47.200 ;
        RECT 145.400 46.200 145.700 46.800 ;
        RECT 146.200 46.200 146.500 46.800 ;
        RECT 145.400 45.800 145.800 46.200 ;
        RECT 146.200 45.800 146.600 46.200 ;
        RECT 139.800 39.800 140.200 40.200 ;
        RECT 132.600 38.800 133.000 39.200 ;
        RECT 132.600 35.200 132.900 38.800 ;
        RECT 139.800 37.200 140.100 39.800 ;
        RECT 135.000 36.800 135.400 37.200 ;
        RECT 136.600 37.100 137.000 37.200 ;
        RECT 137.400 37.100 137.800 37.200 ;
        RECT 136.600 36.800 137.800 37.100 ;
        RECT 139.800 36.800 140.200 37.200 ;
        RECT 135.000 35.200 135.300 36.800 ;
        RECT 135.800 35.800 136.200 36.200 ;
        RECT 135.800 35.200 136.100 35.800 ;
        RECT 132.600 34.800 133.000 35.200 ;
        RECT 133.400 34.800 133.800 35.200 ;
        RECT 135.000 34.800 135.400 35.200 ;
        RECT 135.800 34.800 136.200 35.200 ;
        RECT 133.400 34.200 133.700 34.800 ;
        RECT 133.400 33.800 133.800 34.200 ;
        RECT 136.600 31.800 137.000 32.200 ;
        RECT 140.600 32.100 141.000 37.900 ;
        RECT 142.200 34.800 142.600 35.200 ;
        RECT 142.200 34.200 142.500 34.800 ;
        RECT 142.200 33.800 142.600 34.200 ;
        RECT 143.000 32.800 143.400 33.200 ;
        RECT 127.000 27.100 127.400 27.200 ;
        RECT 127.800 27.100 128.200 27.200 ;
        RECT 126.200 26.800 128.200 27.100 ;
        RECT 131.800 26.800 132.200 27.200 ;
        RECT 132.600 27.100 133.000 27.200 ;
        RECT 133.400 27.100 133.800 27.200 ;
        RECT 132.600 26.800 133.800 27.100 ;
        RECT 131.800 26.200 132.100 26.800 ;
        RECT 119.000 25.800 119.400 26.200 ;
        RECT 119.800 26.100 120.200 26.200 ;
        RECT 120.600 26.100 121.000 26.200 ;
        RECT 119.800 25.800 121.000 26.100 ;
        RECT 121.400 25.800 121.800 26.200 ;
        RECT 123.800 26.100 124.200 26.200 ;
        RECT 124.600 26.100 125.000 26.200 ;
        RECT 123.800 25.800 125.000 26.100 ;
        RECT 126.200 26.100 126.600 26.200 ;
        RECT 127.000 26.100 127.400 26.200 ;
        RECT 126.200 25.800 127.400 26.100 ;
        RECT 131.000 25.800 131.400 26.200 ;
        RECT 131.800 25.800 132.200 26.200 ;
        RECT 116.600 24.800 117.000 25.200 ;
        RECT 119.000 23.200 119.300 25.800 ;
        RECT 119.800 25.100 120.200 25.200 ;
        RECT 120.600 25.100 121.000 25.200 ;
        RECT 119.800 24.800 121.000 25.100 ;
        RECT 124.600 25.100 125.000 25.200 ;
        RECT 125.400 25.100 125.800 25.200 ;
        RECT 124.600 24.800 125.800 25.100 ;
        RECT 129.400 24.800 129.800 25.200 ;
        RECT 118.200 22.800 118.600 23.200 ;
        RECT 119.000 22.800 119.400 23.200 ;
        RECT 118.200 22.200 118.500 22.800 ;
        RECT 118.200 21.800 118.600 22.200 ;
        RECT 129.400 21.200 129.700 24.800 ;
        RECT 130.200 23.800 130.600 24.200 ;
        RECT 115.800 20.800 116.200 21.200 ;
        RECT 129.400 20.800 129.800 21.200 ;
        RECT 130.200 19.200 130.500 23.800 ;
        RECT 130.200 18.800 130.600 19.200 ;
        RECT 115.000 16.800 115.400 17.200 ;
        RECT 115.000 16.100 115.400 16.200 ;
        RECT 115.800 16.100 116.200 16.200 ;
        RECT 113.400 13.100 113.800 15.900 ;
        RECT 115.000 15.800 116.200 16.100 ;
        RECT 117.400 15.800 117.800 16.200 ;
        RECT 115.800 15.200 116.100 15.800 ;
        RECT 117.400 15.200 117.700 15.800 ;
        RECT 115.800 14.800 116.200 15.200 ;
        RECT 117.400 14.800 117.800 15.200 ;
        RECT 118.200 15.100 118.600 15.200 ;
        RECT 119.000 15.100 119.400 15.200 ;
        RECT 118.200 14.800 119.400 15.100 ;
        RECT 114.200 13.800 114.600 14.200 ;
        RECT 118.200 14.100 118.600 14.200 ;
        RECT 119.000 14.100 119.400 14.200 ;
        RECT 118.200 13.800 119.400 14.100 ;
        RECT 114.200 13.200 114.500 13.800 ;
        RECT 114.200 12.800 114.600 13.200 ;
        RECT 119.800 13.100 120.200 15.900 ;
        RECT 120.600 13.800 121.000 14.200 ;
        RECT 120.600 12.200 120.900 13.800 ;
        RECT 120.600 11.800 121.000 12.200 ;
        RECT 121.400 12.100 121.800 17.900 ;
        RECT 122.200 15.800 122.600 16.200 ;
        RECT 122.200 15.100 122.500 15.800 ;
        RECT 122.200 14.700 122.600 15.100 ;
        RECT 125.400 13.800 125.800 14.200 ;
        RECT 125.400 13.200 125.700 13.800 ;
        RECT 125.400 12.800 125.800 13.200 ;
        RECT 126.200 12.100 126.600 17.900 ;
        RECT 107.800 7.800 108.200 8.200 ;
        RECT 105.400 6.800 105.800 7.200 ;
        RECT 108.600 6.800 109.000 7.200 ;
        RECT 105.400 6.200 105.700 6.800 ;
        RECT 108.600 6.300 108.900 6.800 ;
        RECT 105.400 5.800 105.800 6.200 ;
        RECT 108.600 5.900 109.000 6.300 ;
        RECT 109.400 3.100 109.800 8.900 ;
        RECT 110.200 7.200 110.500 11.800 ;
        RECT 131.000 9.200 131.300 25.800 ;
        RECT 135.000 23.100 135.400 28.900 ;
        RECT 136.600 26.200 136.900 31.800 ;
        RECT 142.200 30.800 142.600 31.200 ;
        RECT 136.600 25.800 137.000 26.200 ;
        RECT 139.800 23.100 140.200 28.900 ;
        RECT 142.200 28.200 142.500 30.800 ;
        RECT 143.000 29.200 143.300 32.800 ;
        RECT 145.400 32.100 145.800 37.900 ;
        RECT 146.200 33.800 146.600 34.200 ;
        RECT 143.000 28.800 143.400 29.200 ;
        RECT 144.600 28.800 145.000 29.200 ;
        RECT 144.600 28.200 144.900 28.800 ;
        RECT 140.600 26.800 141.000 27.200 ;
        RECT 140.600 26.200 140.900 26.800 ;
        RECT 140.600 25.800 141.000 26.200 ;
        RECT 136.600 15.800 137.000 16.200 ;
        RECT 136.600 15.200 136.900 15.800 ;
        RECT 136.600 14.800 137.000 15.200 ;
        RECT 137.400 14.800 137.800 15.200 ;
        RECT 137.400 9.200 137.700 14.800 ;
        RECT 139.000 11.800 139.400 12.200 ;
        RECT 111.800 8.800 112.200 9.200 ;
        RECT 119.000 8.800 119.400 9.200 ;
        RECT 122.200 9.100 122.600 9.200 ;
        RECT 123.000 9.100 123.400 9.200 ;
        RECT 122.200 8.800 123.400 9.100 ;
        RECT 110.200 6.800 110.600 7.200 ;
        RECT 111.000 5.100 111.400 7.900 ;
        RECT 111.800 7.200 112.100 8.800 ;
        RECT 119.000 8.200 119.300 8.800 ;
        RECT 116.600 7.800 117.000 8.200 ;
        RECT 119.000 7.800 119.400 8.200 ;
        RECT 121.400 7.800 121.800 8.200 ;
        RECT 116.600 7.200 116.900 7.800 ;
        RECT 121.400 7.200 121.700 7.800 ;
        RECT 111.800 6.800 112.200 7.200 ;
        RECT 113.400 6.800 113.800 7.200 ;
        RECT 116.600 6.800 117.000 7.200 ;
        RECT 117.400 6.800 117.800 7.200 ;
        RECT 121.400 6.800 121.800 7.200 ;
        RECT 113.400 6.200 113.700 6.800 ;
        RECT 116.600 6.200 116.900 6.800 ;
        RECT 117.400 6.200 117.700 6.800 ;
        RECT 113.400 5.800 113.800 6.200 ;
        RECT 115.800 5.800 116.200 6.200 ;
        RECT 116.600 5.800 117.000 6.200 ;
        RECT 117.400 5.800 117.800 6.200 ;
        RECT 120.600 5.800 121.000 6.200 ;
        RECT 121.400 6.100 121.800 6.200 ;
        RECT 122.200 6.100 122.600 6.200 ;
        RECT 121.400 5.800 122.600 6.100 ;
        RECT 115.800 5.200 116.100 5.800 ;
        RECT 120.600 5.200 120.900 5.800 ;
        RECT 112.600 5.100 113.000 5.200 ;
        RECT 113.400 5.100 113.800 5.200 ;
        RECT 112.600 4.800 113.800 5.100 ;
        RECT 115.800 4.800 116.200 5.200 ;
        RECT 120.600 4.800 121.000 5.200 ;
        RECT 125.400 3.100 125.800 8.900 ;
        RECT 127.000 5.800 127.400 6.200 ;
        RECT 127.000 5.200 127.300 5.800 ;
        RECT 127.000 4.800 127.400 5.200 ;
        RECT 130.200 3.100 130.600 8.900 ;
        RECT 131.000 8.800 131.400 9.200 ;
        RECT 132.600 9.100 133.000 9.200 ;
        RECT 133.400 9.100 133.800 9.200 ;
        RECT 132.600 8.800 133.800 9.100 ;
        RECT 131.000 7.800 131.400 8.200 ;
        RECT 131.000 7.200 131.300 7.800 ;
        RECT 131.000 6.800 131.400 7.200 ;
        RECT 131.800 5.100 132.200 7.900 ;
        RECT 136.600 3.100 137.000 8.900 ;
        RECT 137.400 8.800 137.800 9.200 ;
        RECT 137.400 7.800 137.800 8.200 ;
        RECT 137.400 7.200 137.700 7.800 ;
        RECT 137.400 6.800 137.800 7.200 ;
        RECT 139.000 6.200 139.300 11.800 ;
        RECT 140.600 8.200 140.900 25.800 ;
        RECT 141.400 25.100 141.800 27.900 ;
        RECT 142.200 27.800 142.600 28.200 ;
        RECT 144.600 27.800 145.000 28.200 ;
        RECT 146.200 27.200 146.500 33.800 ;
        RECT 147.000 33.100 147.400 35.900 ;
        RECT 146.200 26.800 146.600 27.200 ;
        RECT 143.800 26.100 144.200 26.200 ;
        RECT 144.600 26.100 145.000 26.200 ;
        RECT 143.800 25.800 145.000 26.100 ;
        RECT 146.200 24.200 146.500 26.800 ;
        RECT 146.200 23.800 146.600 24.200 ;
        RECT 147.000 23.100 147.400 28.900 ;
        RECT 147.800 27.200 148.100 46.800 ;
        RECT 148.600 46.200 148.900 46.800 ;
        RECT 159.800 46.200 160.100 46.800 ;
        RECT 148.600 45.800 149.000 46.200 ;
        RECT 151.000 45.800 151.400 46.200 ;
        RECT 155.800 45.800 156.200 46.200 ;
        RECT 157.400 46.100 157.800 46.200 ;
        RECT 156.600 45.800 157.800 46.100 ;
        RECT 159.800 45.800 160.200 46.200 ;
        RECT 148.600 45.100 149.000 45.200 ;
        RECT 149.400 45.100 149.800 45.200 ;
        RECT 148.600 44.800 149.800 45.100 ;
        RECT 151.000 44.200 151.300 45.800 ;
        RECT 155.800 45.200 156.100 45.800 ;
        RECT 155.800 44.800 156.200 45.200 ;
        RECT 151.000 43.800 151.400 44.200 ;
        RECT 148.600 42.800 149.000 43.200 ;
        RECT 148.600 39.200 148.900 42.800 ;
        RECT 155.000 41.800 155.400 42.200 ;
        RECT 148.600 38.800 149.000 39.200 ;
        RECT 154.200 39.100 154.600 39.200 ;
        RECT 155.000 39.100 155.300 41.800 ;
        RECT 154.200 38.800 155.300 39.100 ;
        RECT 151.000 29.800 151.400 30.200 ;
        RECT 147.800 26.800 148.200 27.200 ;
        RECT 151.000 26.300 151.300 29.800 ;
        RECT 148.600 25.800 149.000 26.200 ;
        RECT 151.000 25.900 151.400 26.300 ;
        RECT 142.200 17.800 142.600 18.200 ;
        RECT 146.200 18.100 146.600 18.200 ;
        RECT 147.000 18.100 147.400 18.200 ;
        RECT 146.200 17.800 147.400 18.100 ;
        RECT 141.400 16.800 141.800 17.200 ;
        RECT 141.400 15.200 141.700 16.800 ;
        RECT 141.400 14.800 141.800 15.200 ;
        RECT 142.200 14.100 142.500 17.800 ;
        RECT 148.600 17.200 148.900 25.800 ;
        RECT 151.800 23.100 152.200 28.900 ;
        RECT 153.400 25.100 153.800 27.900 ;
        RECT 154.200 26.200 154.500 38.800 ;
        RECT 155.800 36.200 156.100 44.800 ;
        RECT 156.600 44.200 156.900 45.800 ;
        RECT 156.600 43.800 157.000 44.200 ;
        RECT 156.600 39.200 156.900 43.800 ;
        RECT 159.000 41.800 159.400 42.200 ;
        RECT 156.600 38.800 157.000 39.200 ;
        RECT 159.000 38.200 159.300 41.800 ;
        RECT 160.600 39.200 160.900 67.800 ;
        RECT 162.200 63.100 162.600 68.900 ;
        RECT 163.000 68.200 163.300 73.800 ;
        RECT 163.800 72.800 164.200 73.200 ;
        RECT 163.000 67.800 163.400 68.200 ;
        RECT 163.800 65.200 164.100 72.800 ;
        RECT 163.800 64.800 164.200 65.200 ;
        RECT 163.000 63.800 163.400 64.200 ;
        RECT 164.600 64.100 164.900 85.800 ;
        RECT 165.400 76.200 165.700 87.800 ;
        RECT 166.200 86.100 166.600 86.200 ;
        RECT 167.000 86.100 167.400 86.200 ;
        RECT 166.200 85.800 167.400 86.100 ;
        RECT 167.800 78.200 168.100 91.800 ;
        RECT 168.600 83.100 169.000 88.900 ;
        RECT 170.200 85.100 170.600 87.900 ;
        RECT 171.000 87.200 171.300 93.800 ;
        RECT 171.800 91.800 172.200 92.200 ;
        RECT 171.000 86.800 171.400 87.200 ;
        RECT 171.000 86.200 171.300 86.800 ;
        RECT 171.800 86.200 172.100 91.800 ;
        RECT 171.000 85.800 171.400 86.200 ;
        RECT 171.800 85.800 172.200 86.200 ;
        RECT 171.000 85.100 171.400 85.200 ;
        RECT 171.800 85.100 172.200 85.200 ;
        RECT 171.000 84.800 172.200 85.100 ;
        RECT 172.600 84.200 172.900 94.800 ;
        RECT 173.400 93.200 173.700 104.800 ;
        RECT 179.800 103.100 180.200 108.900 ;
        RECT 180.600 105.200 180.900 121.800 ;
        RECT 188.600 121.200 188.900 121.800 ;
        RECT 191.000 121.200 191.300 121.800 ;
        RECT 188.600 120.800 189.000 121.200 ;
        RECT 191.000 120.800 191.400 121.200 ;
        RECT 183.800 118.800 184.200 119.200 ;
        RECT 183.800 118.200 184.100 118.800 ;
        RECT 183.800 117.800 184.200 118.200 ;
        RECT 185.400 111.800 185.800 112.200 ;
        RECT 187.800 112.100 188.200 117.900 ;
        RECT 188.600 114.800 189.000 115.200 ;
        RECT 191.000 114.800 191.400 115.200 ;
        RECT 188.600 114.200 188.900 114.800 ;
        RECT 191.000 114.200 191.300 114.800 ;
        RECT 188.600 113.800 189.000 114.200 ;
        RECT 191.000 113.800 191.400 114.200 ;
        RECT 185.400 110.200 185.700 111.800 ;
        RECT 185.400 109.800 185.800 110.200 ;
        RECT 183.800 105.900 184.200 106.300 ;
        RECT 183.800 105.200 184.100 105.900 ;
        RECT 180.600 104.800 181.000 105.200 ;
        RECT 183.800 104.800 184.200 105.200 ;
        RECT 182.200 103.800 182.600 104.200 ;
        RECT 182.200 99.200 182.500 103.800 ;
        RECT 184.600 103.100 185.000 108.900 ;
        RECT 185.400 106.800 185.800 107.200 ;
        RECT 182.200 98.800 182.600 99.200 ;
        RECT 179.800 96.100 180.200 96.200 ;
        RECT 180.600 96.100 181.000 96.200 ;
        RECT 179.800 95.800 181.000 96.100 ;
        RECT 182.200 95.200 182.500 98.800 ;
        RECT 185.400 97.200 185.700 106.800 ;
        RECT 186.200 105.100 186.600 107.900 ;
        RECT 187.000 106.800 187.400 107.200 ;
        RECT 187.000 106.200 187.300 106.800 ;
        RECT 191.800 106.200 192.100 125.800 ;
        RECT 192.600 112.100 193.000 117.900 ;
        RECT 194.200 113.100 194.600 115.900 ;
        RECT 195.000 113.100 195.400 115.900 ;
        RECT 196.600 112.100 197.000 117.900 ;
        RECT 197.400 115.100 197.700 126.800 ;
        RECT 198.200 124.200 198.500 126.800 ;
        RECT 199.800 126.100 200.200 126.200 ;
        RECT 200.600 126.100 201.000 126.200 ;
        RECT 199.800 125.800 201.000 126.100 ;
        RECT 198.200 123.800 198.600 124.200 ;
        RECT 197.400 114.700 197.800 115.100 ;
        RECT 198.200 112.200 198.500 123.800 ;
        RECT 203.800 119.200 204.100 126.800 ;
        RECT 204.600 125.800 205.000 126.200 ;
        RECT 204.600 124.200 204.900 125.800 ;
        RECT 204.600 123.800 205.000 124.200 ;
        RECT 203.800 118.800 204.200 119.200 ;
        RECT 199.000 114.800 199.400 115.200 ;
        RECT 198.200 111.800 198.600 112.200 ;
        RECT 196.600 110.800 197.000 111.200 ;
        RECT 192.600 107.800 193.000 108.200 ;
        RECT 192.600 106.200 192.900 107.800 ;
        RECT 196.600 107.200 196.900 110.800 ;
        RECT 199.000 109.200 199.300 114.800 ;
        RECT 201.400 112.100 201.800 117.900 ;
        RECT 202.200 115.800 202.600 116.200 ;
        RECT 201.400 109.800 201.800 110.200 ;
        RECT 199.000 108.800 199.400 109.200 ;
        RECT 201.400 107.200 201.700 109.800 ;
        RECT 196.600 107.100 197.000 107.200 ;
        RECT 197.400 107.100 197.800 107.200 ;
        RECT 196.600 106.800 197.800 107.100 ;
        RECT 199.800 106.800 200.200 107.200 ;
        RECT 201.400 106.800 201.800 107.200 ;
        RECT 187.000 105.800 187.400 106.200 ;
        RECT 187.800 105.800 188.200 106.200 ;
        RECT 190.200 106.100 190.600 106.200 ;
        RECT 191.000 106.100 191.400 106.200 ;
        RECT 190.200 105.800 191.400 106.100 ;
        RECT 191.800 105.800 192.200 106.200 ;
        RECT 192.600 105.800 193.000 106.200 ;
        RECT 195.000 106.100 195.400 106.200 ;
        RECT 195.800 106.100 196.200 106.200 ;
        RECT 195.000 105.800 196.200 106.100 ;
        RECT 196.600 105.800 197.000 106.200 ;
        RECT 187.800 104.200 188.100 105.800 ;
        RECT 187.800 103.800 188.200 104.200 ;
        RECT 190.200 103.200 190.500 105.800 ;
        RECT 190.200 102.800 190.600 103.200 ;
        RECT 189.400 101.800 189.800 102.200 ;
        RECT 185.400 96.800 185.800 97.200 ;
        RECT 176.600 94.800 177.000 95.200 ;
        RECT 177.400 94.800 177.800 95.200 ;
        RECT 178.200 94.800 178.600 95.200 ;
        RECT 180.600 94.800 181.000 95.200 ;
        RECT 182.200 94.800 182.600 95.200 ;
        RECT 175.000 94.100 175.400 94.200 ;
        RECT 175.800 94.100 176.200 94.200 ;
        RECT 175.000 93.800 176.200 94.100 ;
        RECT 173.400 93.100 173.800 93.200 ;
        RECT 174.200 93.100 174.600 93.200 ;
        RECT 173.400 92.800 174.600 93.100 ;
        RECT 174.200 89.800 174.600 90.200 ;
        RECT 174.200 85.200 174.500 89.800 ;
        RECT 176.600 89.200 176.900 94.800 ;
        RECT 177.400 91.200 177.700 94.800 ;
        RECT 178.200 92.200 178.500 94.800 ;
        RECT 178.200 91.800 178.600 92.200 ;
        RECT 177.400 90.800 177.800 91.200 ;
        RECT 178.200 89.800 178.600 90.200 ;
        RECT 175.800 88.800 176.200 89.200 ;
        RECT 176.600 88.800 177.000 89.200 ;
        RECT 175.800 87.200 176.100 88.800 ;
        RECT 175.800 86.800 176.200 87.200 ;
        RECT 178.200 86.200 178.500 89.800 ;
        RECT 179.000 89.100 179.400 89.200 ;
        RECT 179.800 89.100 180.200 89.200 ;
        RECT 179.000 88.800 180.200 89.100 ;
        RECT 179.000 87.800 179.400 88.200 ;
        RECT 179.000 87.200 179.300 87.800 ;
        RECT 179.000 86.800 179.400 87.200 ;
        RECT 176.600 86.100 177.000 86.200 ;
        RECT 177.400 86.100 177.800 86.200 ;
        RECT 176.600 85.800 177.800 86.100 ;
        RECT 178.200 85.800 178.600 86.200 ;
        RECT 173.400 84.800 173.800 85.200 ;
        RECT 174.200 84.800 174.600 85.200 ;
        RECT 171.000 83.800 171.400 84.200 ;
        RECT 172.600 83.800 173.000 84.200 ;
        RECT 171.000 79.200 171.300 83.800 ;
        RECT 171.000 78.800 171.400 79.200 ;
        RECT 167.800 77.800 168.200 78.200 ;
        RECT 172.600 76.800 173.000 77.200 ;
        RECT 165.400 75.800 165.800 76.200 ;
        RECT 167.800 75.800 168.200 76.200 ;
        RECT 165.400 75.200 165.700 75.800 ;
        RECT 165.400 74.800 165.800 75.200 ;
        RECT 167.800 74.200 168.100 75.800 ;
        RECT 168.600 74.800 169.000 75.200 ;
        RECT 169.400 74.800 169.800 75.200 ;
        RECT 167.800 73.800 168.200 74.200 ;
        RECT 168.600 72.200 168.900 74.800 ;
        RECT 169.400 73.200 169.700 74.800 ;
        RECT 172.600 73.200 172.900 76.800 ;
        RECT 173.400 75.200 173.700 84.800 ;
        RECT 175.800 76.800 176.200 77.200 ;
        RECT 175.800 75.200 176.100 76.800 ;
        RECT 180.600 75.200 180.900 94.800 ;
        RECT 186.200 92.100 186.600 97.900 ;
        RECT 189.400 95.200 189.700 101.800 ;
        RECT 190.200 100.800 190.600 101.200 ;
        RECT 189.400 94.800 189.800 95.200 ;
        RECT 189.400 93.800 189.800 94.200 ;
        RECT 182.200 83.100 182.600 88.900 ;
        RECT 183.000 85.800 183.400 86.200 ;
        RECT 184.600 86.100 185.000 86.200 ;
        RECT 185.400 86.100 185.800 86.200 ;
        RECT 184.600 85.800 185.800 86.100 ;
        RECT 183.000 77.200 183.300 85.800 ;
        RECT 185.400 84.800 185.800 85.200 ;
        RECT 181.400 76.800 181.800 77.200 ;
        RECT 183.000 76.800 183.400 77.200 ;
        RECT 181.400 76.200 181.700 76.800 ;
        RECT 181.400 75.800 181.800 76.200 ;
        RECT 173.400 74.800 173.800 75.200 ;
        RECT 175.800 74.800 176.200 75.200 ;
        RECT 176.600 75.100 177.000 75.200 ;
        RECT 177.400 75.100 177.800 75.200 ;
        RECT 176.600 74.800 177.800 75.100 ;
        RECT 179.800 74.800 180.200 75.200 ;
        RECT 180.600 74.800 181.000 75.200 ;
        RECT 173.400 74.100 173.800 74.200 ;
        RECT 174.200 74.100 174.600 74.200 ;
        RECT 173.400 73.800 174.600 74.100 ;
        RECT 175.800 73.200 176.100 74.800 ;
        RECT 179.800 74.200 180.100 74.800 ;
        RECT 178.200 74.100 178.600 74.200 ;
        RECT 179.000 74.100 179.400 74.200 ;
        RECT 178.200 73.800 179.400 74.100 ;
        RECT 179.800 73.800 180.200 74.200 ;
        RECT 169.400 72.800 169.800 73.200 ;
        RECT 172.600 72.800 173.000 73.200 ;
        RECT 175.800 72.800 176.200 73.200 ;
        RECT 167.000 71.800 167.400 72.200 ;
        RECT 168.600 71.800 169.000 72.200 ;
        RECT 165.400 66.800 165.800 67.200 ;
        RECT 166.200 66.800 166.600 67.200 ;
        RECT 165.400 66.200 165.700 66.800 ;
        RECT 166.200 66.200 166.500 66.800 ;
        RECT 165.400 65.800 165.800 66.200 ;
        RECT 166.200 65.800 166.600 66.200 ;
        RECT 165.400 64.100 165.800 64.200 ;
        RECT 164.600 63.800 165.800 64.100 ;
        RECT 162.200 52.100 162.600 57.900 ;
        RECT 163.000 49.200 163.300 63.800 ;
        RECT 165.400 54.200 165.700 63.800 ;
        RECT 167.000 59.200 167.300 71.800 ;
        RECT 180.600 70.200 180.900 74.800 ;
        RECT 183.800 72.100 184.200 77.900 ;
        RECT 184.600 74.800 185.000 75.200 ;
        RECT 184.600 71.200 184.900 74.800 ;
        RECT 181.400 70.800 181.800 71.200 ;
        RECT 184.600 70.800 185.000 71.200 ;
        RECT 180.600 69.800 181.000 70.200 ;
        RECT 169.400 66.800 169.800 67.200 ;
        RECT 169.400 66.200 169.700 66.800 ;
        RECT 167.800 66.100 168.200 66.200 ;
        RECT 168.600 66.100 169.000 66.200 ;
        RECT 167.800 65.800 169.000 66.100 ;
        RECT 169.400 65.800 169.800 66.200 ;
        RECT 173.400 65.800 173.800 66.200 ;
        RECT 167.800 65.100 168.200 65.200 ;
        RECT 168.600 65.100 169.000 65.200 ;
        RECT 167.800 64.800 169.000 65.100 ;
        RECT 167.000 58.800 167.400 59.200 ;
        RECT 166.200 54.700 166.600 55.100 ;
        RECT 165.400 53.800 165.800 54.200 ;
        RECT 161.400 48.800 161.800 49.200 ;
        RECT 163.000 48.800 163.400 49.200 ;
        RECT 161.400 46.200 161.700 48.800 ;
        RECT 162.200 46.800 162.600 47.200 ;
        RECT 161.400 45.800 161.800 46.200 ;
        RECT 162.200 40.200 162.500 46.800 ;
        RECT 164.600 45.800 165.000 46.200 ;
        RECT 164.600 45.200 164.900 45.800 ;
        RECT 164.600 44.800 165.000 45.200 ;
        RECT 164.600 43.800 165.000 44.200 ;
        RECT 162.200 39.800 162.600 40.200 ;
        RECT 160.600 38.800 161.000 39.200 ;
        RECT 163.000 38.800 163.400 39.200 ;
        RECT 159.000 37.800 159.400 38.200 ;
        RECT 155.800 35.800 156.200 36.200 ;
        RECT 160.600 32.100 161.000 37.900 ;
        RECT 162.200 37.800 162.600 38.200 ;
        RECT 162.200 35.200 162.500 37.800 ;
        RECT 162.200 34.800 162.600 35.200 ;
        RECT 161.400 30.800 161.800 31.200 ;
        RECT 157.400 29.800 157.800 30.200 ;
        RECT 157.400 29.200 157.700 29.800 ;
        RECT 157.400 28.800 157.800 29.200 ;
        RECT 161.400 28.200 161.700 30.800 ;
        RECT 163.000 28.200 163.300 38.800 ;
        RECT 164.600 29.200 164.900 43.800 ;
        RECT 165.400 43.200 165.700 53.800 ;
        RECT 166.200 53.200 166.500 54.700 ;
        RECT 166.200 52.800 166.600 53.200 ;
        RECT 167.000 52.100 167.400 57.900 ;
        RECT 168.600 53.100 169.000 55.900 ;
        RECT 169.400 55.800 169.800 56.200 ;
        RECT 169.400 55.200 169.700 55.800 ;
        RECT 173.400 55.200 173.700 65.800 ;
        RECT 174.200 63.100 174.600 68.900 ;
        RECT 175.000 65.800 175.400 66.200 ;
        RECT 175.800 65.800 176.200 66.200 ;
        RECT 175.000 64.200 175.300 65.800 ;
        RECT 175.800 65.200 176.100 65.800 ;
        RECT 175.800 64.800 176.200 65.200 ;
        RECT 177.400 64.800 177.800 65.200 ;
        RECT 175.000 63.800 175.400 64.200 ;
        RECT 176.600 61.800 177.000 62.200 ;
        RECT 176.600 59.200 176.900 61.800 ;
        RECT 176.600 58.800 177.000 59.200 ;
        RECT 177.400 56.200 177.700 64.800 ;
        RECT 179.000 63.100 179.400 68.900 ;
        RECT 180.600 65.100 181.000 67.900 ;
        RECT 181.400 67.200 181.700 70.800 ;
        RECT 182.200 69.800 182.600 70.200 ;
        RECT 181.400 66.800 181.800 67.200 ;
        RECT 182.200 66.200 182.500 69.800 ;
        RECT 185.400 66.200 185.700 84.800 ;
        RECT 187.000 83.100 187.400 88.900 ;
        RECT 188.600 85.100 189.000 87.900 ;
        RECT 189.400 87.200 189.700 93.800 ;
        RECT 189.400 86.800 189.800 87.200 ;
        RECT 190.200 86.200 190.500 100.800 ;
        RECT 191.000 92.100 191.400 97.900 ;
        RECT 191.000 86.800 191.400 87.200 ;
        RECT 191.000 86.200 191.300 86.800 ;
        RECT 190.200 85.800 190.600 86.200 ;
        RECT 191.000 85.800 191.400 86.200 ;
        RECT 190.200 83.200 190.500 85.800 ;
        RECT 191.800 85.200 192.100 105.800 ;
        RECT 194.200 105.100 194.600 105.200 ;
        RECT 195.000 105.100 195.400 105.200 ;
        RECT 194.200 104.800 195.400 105.100 ;
        RECT 192.600 93.100 193.000 95.900 ;
        RECT 192.600 92.100 193.000 92.200 ;
        RECT 193.400 92.100 193.800 92.200 ;
        RECT 192.600 91.800 193.800 92.100 ;
        RECT 196.600 88.200 196.900 105.800 ;
        RECT 199.800 105.200 200.100 106.800 ;
        RECT 202.200 105.200 202.500 115.800 ;
        RECT 199.800 104.800 200.200 105.200 ;
        RECT 202.200 104.800 202.600 105.200 ;
        RECT 202.200 103.200 202.500 104.800 ;
        RECT 202.200 102.800 202.600 103.200 ;
        RECT 202.200 102.100 202.600 102.200 ;
        RECT 203.000 102.100 203.400 102.200 ;
        RECT 202.200 101.800 203.400 102.100 ;
        RECT 197.400 92.100 197.800 97.900 ;
        RECT 200.600 95.800 201.000 96.200 ;
        RECT 200.600 95.200 200.900 95.800 ;
        RECT 198.200 94.800 198.600 95.200 ;
        RECT 200.600 94.800 201.000 95.200 ;
        RECT 198.200 94.200 198.500 94.800 ;
        RECT 198.200 93.800 198.600 94.200 ;
        RECT 201.400 92.800 201.800 93.200 ;
        RECT 196.600 87.800 197.000 88.200 ;
        RECT 192.600 86.800 193.000 87.200 ;
        RECT 192.600 86.200 192.900 86.800 ;
        RECT 192.600 85.800 193.000 86.200 ;
        RECT 193.400 85.800 193.800 86.200 ;
        RECT 194.200 86.100 194.600 86.200 ;
        RECT 195.000 86.100 195.400 86.200 ;
        RECT 194.200 85.800 195.400 86.100 ;
        RECT 193.400 85.200 193.700 85.800 ;
        RECT 191.800 84.800 192.200 85.200 ;
        RECT 193.400 84.800 193.800 85.200 ;
        RECT 191.000 83.800 191.400 84.200 ;
        RECT 190.200 82.800 190.600 83.200 ;
        RECT 191.000 79.200 191.300 83.800 ;
        RECT 191.000 78.800 191.400 79.200 ;
        RECT 186.200 74.800 186.600 75.200 ;
        RECT 186.200 74.200 186.500 74.800 ;
        RECT 186.200 73.800 186.600 74.200 ;
        RECT 188.600 72.100 189.000 77.900 ;
        RECT 190.200 73.100 190.600 75.900 ;
        RECT 192.600 74.800 193.000 75.200 ;
        RECT 195.000 75.100 195.400 75.200 ;
        RECT 195.800 75.100 196.200 75.200 ;
        RECT 195.000 74.800 196.200 75.100 ;
        RECT 191.800 73.800 192.200 74.200 ;
        RECT 191.800 73.200 192.100 73.800 ;
        RECT 191.800 72.800 192.200 73.200 ;
        RECT 192.600 73.100 192.900 74.800 ;
        RECT 193.400 74.100 193.800 74.200 ;
        RECT 194.200 74.100 194.600 74.200 ;
        RECT 193.400 73.800 194.600 74.100 ;
        RECT 192.600 72.800 193.700 73.100 ;
        RECT 187.000 69.800 187.400 70.200 ;
        RECT 187.000 67.200 187.300 69.800 ;
        RECT 193.400 69.200 193.700 72.800 ;
        RECT 187.800 68.800 188.200 69.200 ;
        RECT 193.400 68.800 193.800 69.200 ;
        RECT 187.800 68.200 188.100 68.800 ;
        RECT 187.800 67.800 188.200 68.200 ;
        RECT 186.200 66.800 186.600 67.200 ;
        RECT 187.000 66.800 187.400 67.200 ;
        RECT 191.000 67.100 191.400 67.200 ;
        RECT 191.800 67.100 192.200 67.200 ;
        RECT 191.000 66.800 192.200 67.100 ;
        RECT 186.200 66.200 186.500 66.800 ;
        RECT 182.200 65.800 182.600 66.200 ;
        RECT 184.600 65.800 185.000 66.200 ;
        RECT 185.400 65.800 185.800 66.200 ;
        RECT 186.200 65.800 186.600 66.200 ;
        RECT 191.000 65.800 191.400 66.200 ;
        RECT 191.800 65.800 192.200 66.200 ;
        RECT 184.600 64.200 184.900 65.800 ;
        RECT 184.600 63.800 185.000 64.200 ;
        RECT 183.000 61.800 183.400 62.200 ;
        RECT 177.400 55.800 177.800 56.200 ;
        RECT 169.400 54.800 169.800 55.200 ;
        RECT 170.200 54.800 170.600 55.200 ;
        RECT 173.400 54.800 173.800 55.200 ;
        RECT 174.200 54.800 174.600 55.200 ;
        RECT 170.200 54.200 170.500 54.800 ;
        RECT 170.200 53.800 170.600 54.200 ;
        RECT 171.000 53.100 171.400 53.200 ;
        RECT 171.800 53.100 172.200 53.200 ;
        RECT 171.000 52.800 172.200 53.100 ;
        RECT 174.200 51.200 174.500 54.800 ;
        RECT 175.000 53.800 175.400 54.200 ;
        RECT 175.000 53.200 175.300 53.800 ;
        RECT 175.000 52.800 175.400 53.200 ;
        RECT 167.000 50.800 167.400 51.200 ;
        RECT 174.200 50.800 174.600 51.200 ;
        RECT 167.000 49.200 167.300 50.800 ;
        RECT 170.200 49.800 170.600 50.200 ;
        RECT 167.000 48.800 167.400 49.200 ;
        RECT 167.000 47.200 167.300 48.800 ;
        RECT 167.000 46.800 167.400 47.200 ;
        RECT 167.000 45.800 167.400 46.200 ;
        RECT 165.400 42.800 165.800 43.200 ;
        RECT 167.000 39.200 167.300 45.800 ;
        RECT 170.200 45.200 170.500 49.800 ;
        RECT 170.200 44.800 170.600 45.200 ;
        RECT 175.000 45.100 175.400 47.900 ;
        RECT 176.600 43.100 177.000 48.900 ;
        RECT 177.400 46.200 177.700 55.800 ;
        RECT 179.000 54.800 179.400 55.200 ;
        RECT 179.800 54.800 180.200 55.200 ;
        RECT 179.000 54.200 179.300 54.800 ;
        RECT 179.800 54.200 180.100 54.800 ;
        RECT 179.000 53.800 179.400 54.200 ;
        RECT 179.800 53.800 180.200 54.200 ;
        RECT 180.600 53.100 181.000 55.900 ;
        RECT 181.400 53.800 181.800 54.200 ;
        RECT 181.400 52.100 181.700 53.800 ;
        RECT 182.200 52.100 182.600 57.900 ;
        RECT 183.000 55.100 183.300 61.800 ;
        RECT 183.000 54.700 183.400 55.100 ;
        RECT 184.600 53.800 185.000 54.200 ;
        RECT 185.400 54.100 185.700 65.800 ;
        RECT 186.200 55.200 186.500 65.800 ;
        RECT 188.600 65.100 189.000 65.200 ;
        RECT 189.400 65.100 189.800 65.200 ;
        RECT 188.600 64.800 189.800 65.100 ;
        RECT 189.400 62.200 189.700 64.800 ;
        RECT 191.000 64.200 191.300 65.800 ;
        RECT 191.800 65.200 192.100 65.800 ;
        RECT 191.800 64.800 192.200 65.200 ;
        RECT 191.000 63.800 191.400 64.200 ;
        RECT 189.400 61.800 189.800 62.200 ;
        RECT 191.000 59.200 191.300 63.800 ;
        RECT 192.600 62.800 193.000 63.200 ;
        RECT 192.600 59.200 192.900 62.800 ;
        RECT 191.000 58.800 191.400 59.200 ;
        RECT 192.600 58.800 193.000 59.200 ;
        RECT 186.200 54.800 186.600 55.200 ;
        RECT 185.400 53.800 186.500 54.100 ;
        RECT 180.600 51.800 181.700 52.100 ;
        RECT 178.200 47.800 178.600 48.200 ;
        RECT 178.200 46.200 178.500 47.800 ;
        RECT 180.600 46.200 180.900 51.800 ;
        RECT 177.400 45.800 177.800 46.200 ;
        RECT 178.200 45.800 178.600 46.200 ;
        RECT 180.600 45.800 181.000 46.200 ;
        RECT 167.800 42.100 168.200 42.200 ;
        RECT 168.600 42.100 169.000 42.200 ;
        RECT 167.800 41.800 169.000 42.100 ;
        RECT 170.200 42.100 170.600 42.200 ;
        RECT 171.000 42.100 171.400 42.200 ;
        RECT 170.200 41.800 171.400 42.100 ;
        RECT 173.400 42.100 173.800 42.200 ;
        RECT 174.200 42.100 174.600 42.200 ;
        RECT 173.400 41.800 174.600 42.100 ;
        RECT 173.400 41.200 173.700 41.800 ;
        RECT 173.400 40.800 173.800 41.200 ;
        RECT 167.800 39.800 168.200 40.200 ;
        RECT 167.000 38.800 167.400 39.200 ;
        RECT 165.400 32.100 165.800 37.900 ;
        RECT 166.200 33.800 166.600 34.200 ;
        RECT 166.200 33.200 166.500 33.800 ;
        RECT 166.200 32.800 166.600 33.200 ;
        RECT 167.000 33.100 167.400 35.900 ;
        RECT 167.800 33.200 168.100 39.800 ;
        RECT 169.400 37.800 169.800 38.200 ;
        RECT 171.800 37.800 172.200 38.200 ;
        RECT 169.400 35.200 169.700 37.800 ;
        RECT 169.400 34.800 169.800 35.200 ;
        RECT 171.800 34.200 172.100 37.800 ;
        RECT 173.400 36.800 173.800 37.200 ;
        RECT 173.400 35.200 173.700 36.800 ;
        RECT 174.200 35.800 174.600 36.200 ;
        RECT 178.200 36.100 178.600 36.200 ;
        RECT 179.000 36.100 179.400 36.200 ;
        RECT 178.200 35.800 179.400 36.100 ;
        RECT 174.200 35.200 174.500 35.800 ;
        RECT 180.600 35.200 180.900 45.800 ;
        RECT 181.400 43.100 181.800 48.900 ;
        RECT 184.600 46.200 184.900 53.800 ;
        RECT 186.200 46.200 186.500 53.800 ;
        RECT 187.000 52.100 187.400 57.900 ;
        RECT 191.800 56.100 192.200 56.200 ;
        RECT 192.600 56.100 193.000 56.200 ;
        RECT 191.800 55.800 193.000 56.100 ;
        RECT 190.200 54.800 190.600 55.200 ;
        RECT 187.800 48.100 188.200 48.200 ;
        RECT 188.600 48.100 189.000 48.200 ;
        RECT 187.800 47.800 189.000 48.100 ;
        RECT 190.200 47.200 190.500 54.800 ;
        RECT 191.800 50.200 192.100 55.800 ;
        RECT 194.200 55.200 194.500 73.800 ;
        RECT 195.000 73.100 195.400 73.200 ;
        RECT 195.800 73.100 196.200 73.200 ;
        RECT 195.000 72.800 196.200 73.100 ;
        RECT 195.000 68.800 195.400 69.200 ;
        RECT 195.000 68.200 195.300 68.800 ;
        RECT 196.600 68.200 196.900 87.800 ;
        RECT 198.200 83.100 198.600 88.900 ;
        RECT 201.400 87.200 201.700 92.800 ;
        RECT 202.200 92.100 202.600 97.900 ;
        RECT 203.800 93.100 204.200 95.900 ;
        RECT 201.400 86.800 201.800 87.200 ;
        RECT 202.200 86.800 202.600 87.200 ;
        RECT 200.600 86.100 201.000 86.200 ;
        RECT 201.400 86.100 201.800 86.200 ;
        RECT 200.600 85.800 201.800 86.100 ;
        RECT 197.400 72.800 197.800 73.200 ;
        RECT 197.400 70.200 197.700 72.800 ;
        RECT 198.200 72.100 198.600 77.900 ;
        RECT 199.800 75.100 200.200 75.200 ;
        RECT 200.600 75.100 201.000 75.200 ;
        RECT 199.800 74.800 201.000 75.100 ;
        RECT 202.200 74.200 202.500 86.800 ;
        RECT 203.000 83.100 203.400 88.900 ;
        RECT 204.600 85.100 205.000 87.900 ;
        RECT 203.800 82.800 204.200 83.200 ;
        RECT 199.800 73.800 200.200 74.200 ;
        RECT 202.200 73.800 202.600 74.200 ;
        RECT 199.000 72.800 199.400 73.200 ;
        RECT 197.400 69.800 197.800 70.200 ;
        RECT 195.000 67.800 195.400 68.200 ;
        RECT 196.600 67.800 197.000 68.200 ;
        RECT 197.400 68.100 197.700 69.800 ;
        RECT 199.000 69.200 199.300 72.800 ;
        RECT 199.000 68.800 199.400 69.200 ;
        RECT 198.200 68.100 198.600 68.200 ;
        RECT 197.400 67.800 198.600 68.100 ;
        RECT 199.000 67.800 199.400 68.200 ;
        RECT 196.600 67.100 197.000 67.200 ;
        RECT 197.400 67.100 197.800 67.200 ;
        RECT 196.600 66.800 197.800 67.100 ;
        RECT 195.800 66.100 196.200 66.200 ;
        RECT 196.600 66.100 197.000 66.200 ;
        RECT 195.800 65.800 197.000 66.100 ;
        RECT 195.000 64.800 195.400 65.200 ;
        RECT 195.000 62.200 195.300 64.800 ;
        RECT 195.000 61.800 195.400 62.200 ;
        RECT 199.000 55.200 199.300 67.800 ;
        RECT 199.800 66.200 200.100 73.800 ;
        RECT 203.000 72.100 203.400 77.900 ;
        RECT 200.600 68.800 201.000 69.200 ;
        RECT 201.400 68.800 201.800 69.200 ;
        RECT 200.600 68.200 200.900 68.800 ;
        RECT 201.400 68.200 201.700 68.800 ;
        RECT 200.600 67.800 201.000 68.200 ;
        RECT 201.400 67.800 201.800 68.200 ;
        RECT 202.200 66.800 202.600 67.200 ;
        RECT 203.000 66.800 203.400 67.200 ;
        RECT 202.200 66.200 202.500 66.800 ;
        RECT 203.000 66.200 203.300 66.800 ;
        RECT 199.800 65.800 200.200 66.200 ;
        RECT 202.200 65.800 202.600 66.200 ;
        RECT 203.000 65.800 203.400 66.200 ;
        RECT 199.800 56.100 200.200 56.200 ;
        RECT 200.600 56.100 201.000 56.200 ;
        RECT 199.800 55.800 201.000 56.100 ;
        RECT 203.800 56.100 204.100 82.800 ;
        RECT 204.600 73.100 205.000 75.900 ;
        RECT 203.800 55.800 204.900 56.100 ;
        RECT 204.600 55.200 204.900 55.800 ;
        RECT 192.600 55.100 193.000 55.200 ;
        RECT 193.400 55.100 193.800 55.200 ;
        RECT 192.600 54.800 193.800 55.100 ;
        RECT 194.200 54.800 194.600 55.200 ;
        RECT 196.600 55.100 197.000 55.200 ;
        RECT 197.400 55.100 197.800 55.200 ;
        RECT 196.600 54.800 197.800 55.100 ;
        RECT 199.000 54.800 199.400 55.200 ;
        RECT 203.800 54.800 204.200 55.200 ;
        RECT 204.600 54.800 205.000 55.200 ;
        RECT 194.200 54.200 194.500 54.800 ;
        RECT 203.800 54.200 204.100 54.800 ;
        RECT 194.200 53.800 194.600 54.200 ;
        RECT 203.800 54.100 204.200 54.200 ;
        RECT 203.800 53.800 204.900 54.100 ;
        RECT 191.800 49.800 192.200 50.200 ;
        RECT 190.200 46.800 190.600 47.200 ;
        RECT 190.200 46.200 190.500 46.800 ;
        RECT 184.600 46.100 185.000 46.200 ;
        RECT 185.400 46.100 185.800 46.200 ;
        RECT 184.600 45.800 185.800 46.100 ;
        RECT 186.200 45.800 186.600 46.200 ;
        RECT 187.000 46.100 187.400 46.200 ;
        RECT 187.800 46.100 188.200 46.200 ;
        RECT 187.000 45.800 188.200 46.100 ;
        RECT 190.200 45.800 190.600 46.200 ;
        RECT 186.200 42.200 186.500 45.800 ;
        RECT 191.000 45.100 191.400 47.900 ;
        RECT 191.800 46.800 192.200 47.200 ;
        RECT 191.800 43.200 192.100 46.800 ;
        RECT 191.800 42.800 192.200 43.200 ;
        RECT 192.600 43.100 193.000 48.900 ;
        RECT 184.600 41.800 185.000 42.200 ;
        RECT 186.200 41.800 186.600 42.200 ;
        RECT 191.800 41.800 192.200 42.200 ;
        RECT 181.400 36.800 181.800 37.200 ;
        RECT 183.800 36.800 184.200 37.200 ;
        RECT 181.400 35.200 181.700 36.800 ;
        RECT 172.600 34.800 173.000 35.200 ;
        RECT 173.400 34.800 173.800 35.200 ;
        RECT 174.200 34.800 174.600 35.200 ;
        RECT 176.600 34.800 177.000 35.200 ;
        RECT 177.400 34.800 177.800 35.200 ;
        RECT 180.600 34.800 181.000 35.200 ;
        RECT 181.400 34.800 181.800 35.200 ;
        RECT 169.400 33.800 169.800 34.200 ;
        RECT 171.800 33.800 172.200 34.200 ;
        RECT 167.800 32.800 168.200 33.200 ;
        RECT 167.800 29.200 168.100 32.800 ;
        RECT 164.600 28.800 165.000 29.200 ;
        RECT 167.800 28.800 168.200 29.200 ;
        RECT 159.000 28.100 159.400 28.200 ;
        RECT 159.800 28.100 160.200 28.200 ;
        RECT 159.000 27.800 160.200 28.100 ;
        RECT 161.400 27.800 161.800 28.200 ;
        RECT 163.000 27.800 163.400 28.200 ;
        RECT 167.000 27.800 167.400 28.200 ;
        RECT 167.800 27.800 168.200 28.200 ;
        RECT 163.000 27.200 163.300 27.800 ;
        RECT 167.000 27.200 167.300 27.800 ;
        RECT 155.800 27.100 156.200 27.200 ;
        RECT 156.600 27.100 157.000 27.200 ;
        RECT 155.800 26.800 157.000 27.100 ;
        RECT 160.600 26.800 161.000 27.200 ;
        RECT 163.000 26.800 163.400 27.200 ;
        RECT 167.000 26.800 167.400 27.200 ;
        RECT 160.600 26.200 160.900 26.800 ;
        RECT 154.200 25.800 154.600 26.200 ;
        RECT 155.800 25.800 156.200 26.200 ;
        RECT 156.600 25.800 157.000 26.200 ;
        RECT 160.600 25.800 161.000 26.200 ;
        RECT 162.200 25.800 162.600 26.200 ;
        RECT 163.800 26.100 164.200 26.200 ;
        RECT 164.600 26.100 165.000 26.200 ;
        RECT 163.800 25.800 165.000 26.100 ;
        RECT 167.000 26.100 167.400 26.200 ;
        RECT 167.800 26.100 168.100 27.800 ;
        RECT 167.000 25.800 168.100 26.100 ;
        RECT 146.200 16.800 146.600 17.200 ;
        RECT 148.600 16.800 149.000 17.200 ;
        RECT 146.200 15.200 146.500 16.800 ;
        RECT 141.400 13.800 142.500 14.100 ;
        RECT 143.000 14.800 143.400 15.200 ;
        RECT 146.200 14.800 146.600 15.200 ;
        RECT 143.000 14.200 143.300 14.800 ;
        RECT 143.000 13.800 143.400 14.200 ;
        RECT 145.400 14.100 145.800 14.200 ;
        RECT 146.200 14.100 146.600 14.200 ;
        RECT 145.400 13.800 146.600 14.100 ;
        RECT 141.400 13.200 141.700 13.800 ;
        RECT 141.400 12.800 141.800 13.200 ;
        RECT 144.600 12.800 145.000 13.200 ;
        RECT 144.600 12.200 144.900 12.800 ;
        RECT 144.600 11.800 145.000 12.200 ;
        RECT 149.400 12.100 149.800 17.900 ;
        RECT 150.200 14.800 150.600 15.200 ;
        RECT 151.000 14.800 151.400 15.200 ;
        RECT 140.600 7.800 141.000 8.200 ;
        RECT 139.000 5.800 139.400 6.200 ;
        RECT 141.400 3.100 141.800 8.900 ;
        RECT 143.000 5.100 143.400 7.900 ;
        RECT 150.200 7.200 150.500 14.800 ;
        RECT 151.000 13.200 151.300 14.800 ;
        RECT 151.000 12.800 151.400 13.200 ;
        RECT 154.200 12.100 154.600 17.900 ;
        RECT 155.800 17.200 156.100 25.800 ;
        RECT 155.800 16.800 156.200 17.200 ;
        RECT 155.800 13.100 156.200 15.900 ;
        RECT 156.600 13.200 156.900 25.800 ;
        RECT 162.200 25.200 162.500 25.800 ;
        RECT 162.200 24.800 162.600 25.200 ;
        RECT 163.800 25.100 164.200 25.200 ;
        RECT 164.600 25.100 165.000 25.200 ;
        RECT 163.800 24.800 165.000 25.100 ;
        RECT 167.800 24.800 168.200 25.200 ;
        RECT 163.800 18.800 164.200 19.200 ;
        RECT 159.800 17.800 160.200 18.200 ;
        RECT 162.200 17.800 162.600 18.200 ;
        RECT 159.800 15.200 160.100 17.800 ;
        RECT 159.800 14.800 160.200 15.200 ;
        RECT 159.800 14.200 160.100 14.800 ;
        RECT 162.200 14.200 162.500 17.800 ;
        RECT 163.000 16.800 163.400 17.200 ;
        RECT 163.000 15.200 163.300 16.800 ;
        RECT 163.000 14.800 163.400 15.200 ;
        RECT 159.800 13.800 160.200 14.200 ;
        RECT 162.200 13.800 162.600 14.200 ;
        RECT 163.800 13.200 164.100 18.800 ;
        RECT 165.400 15.800 165.800 16.200 ;
        RECT 165.400 15.200 165.700 15.800 ;
        RECT 165.400 14.800 165.800 15.200 ;
        RECT 165.400 14.200 165.700 14.800 ;
        RECT 167.800 14.200 168.100 24.800 ;
        RECT 169.400 24.200 169.700 33.800 ;
        RECT 172.600 32.200 172.900 34.800 ;
        RECT 171.000 32.100 171.400 32.200 ;
        RECT 171.000 31.800 172.100 32.100 ;
        RECT 172.600 31.800 173.000 32.200 ;
        RECT 169.400 23.800 169.800 24.200 ;
        RECT 170.200 23.100 170.600 28.900 ;
        RECT 171.800 26.200 172.100 31.800 ;
        RECT 171.800 25.800 172.200 26.200 ;
        RECT 168.600 16.800 169.000 17.200 ;
        RECT 168.600 15.200 168.900 16.800 ;
        RECT 173.400 15.200 173.700 34.800 ;
        RECT 176.600 32.200 176.900 34.800 ;
        RECT 177.400 34.200 177.700 34.800 ;
        RECT 177.400 33.800 177.800 34.200 ;
        RECT 179.000 33.800 179.400 34.200 ;
        RECT 179.000 33.200 179.300 33.800 ;
        RECT 179.000 32.800 179.400 33.200 ;
        RECT 179.800 32.800 180.200 33.200 ;
        RECT 176.600 31.800 177.000 32.200 ;
        RECT 179.800 32.100 180.100 32.800 ;
        RECT 179.000 31.800 180.100 32.100 ;
        RECT 179.000 29.200 179.300 31.800 ;
        RECT 175.000 23.100 175.400 28.900 ;
        RECT 179.000 28.800 179.400 29.200 ;
        RECT 179.000 28.200 179.300 28.800 ;
        RECT 175.800 26.800 176.200 27.200 ;
        RECT 175.800 26.200 176.100 26.800 ;
        RECT 175.800 25.800 176.200 26.200 ;
        RECT 175.800 15.200 176.100 25.800 ;
        RECT 176.600 25.100 177.000 27.900 ;
        RECT 179.000 27.800 179.400 28.200 ;
        RECT 179.800 23.100 180.200 28.900 ;
        RECT 180.600 27.200 180.900 34.800 ;
        RECT 183.800 34.200 184.100 36.800 ;
        RECT 184.600 35.200 184.900 41.800 ;
        RECT 184.600 35.100 185.000 35.200 ;
        RECT 184.600 34.800 185.700 35.100 ;
        RECT 183.800 33.800 184.200 34.200 ;
        RECT 184.600 33.800 185.000 34.200 ;
        RECT 184.600 33.200 184.900 33.800 ;
        RECT 184.600 32.800 185.000 33.200 ;
        RECT 181.400 31.800 181.800 32.200 ;
        RECT 183.000 31.800 183.400 32.200 ;
        RECT 181.400 27.200 181.700 31.800 ;
        RECT 180.600 26.800 181.000 27.200 ;
        RECT 181.400 26.800 181.800 27.200 ;
        RECT 180.600 26.200 180.900 26.800 ;
        RECT 180.600 25.800 181.000 26.200 ;
        RECT 178.200 17.800 178.600 18.200 ;
        RECT 180.600 17.800 181.000 18.200 ;
        RECT 178.200 15.200 178.500 17.800 ;
        RECT 168.600 14.800 169.000 15.200 ;
        RECT 173.400 14.800 173.800 15.200 ;
        RECT 175.800 14.800 176.200 15.200 ;
        RECT 178.200 14.800 178.600 15.200 ;
        RECT 165.400 13.800 165.800 14.200 ;
        RECT 167.800 13.800 168.200 14.200 ;
        RECT 156.600 12.800 157.000 13.200 ;
        RECT 163.000 12.800 163.400 13.200 ;
        RECT 163.800 12.800 164.200 13.200 ;
        RECT 156.600 9.200 156.900 12.800 ;
        RECT 161.400 11.800 161.800 12.200 ;
        RECT 161.400 9.200 161.700 11.800 ;
        RECT 162.200 9.800 162.600 10.200 ;
        RECT 152.600 9.100 153.000 9.200 ;
        RECT 153.400 9.100 153.800 9.200 ;
        RECT 152.600 8.800 153.800 9.100 ;
        RECT 150.200 6.800 150.600 7.200 ;
        RECT 155.000 3.100 155.400 8.900 ;
        RECT 156.600 8.800 157.000 9.200 ;
        RECT 159.000 8.800 159.400 9.200 ;
        RECT 159.000 6.300 159.300 8.800 ;
        RECT 159.000 5.900 159.400 6.300 ;
        RECT 159.800 3.100 160.200 8.900 ;
        RECT 161.400 8.800 161.800 9.200 ;
        RECT 162.200 8.200 162.500 9.800 ;
        RECT 163.000 9.200 163.300 12.800 ;
        RECT 163.800 9.200 164.100 12.800 ;
        RECT 167.000 11.800 167.400 12.200 ;
        RECT 163.000 8.800 163.400 9.200 ;
        RECT 163.800 8.800 164.200 9.200 ;
        RECT 160.600 7.800 161.000 8.200 ;
        RECT 160.600 7.200 160.900 7.800 ;
        RECT 160.600 6.800 161.000 7.200 ;
        RECT 161.400 5.100 161.800 7.900 ;
        RECT 162.200 7.800 162.600 8.200 ;
        RECT 166.200 3.100 166.600 8.900 ;
        RECT 167.000 6.100 167.300 11.800 ;
        RECT 173.400 10.800 173.800 11.200 ;
        RECT 173.400 9.200 173.700 10.800 ;
        RECT 175.800 10.100 176.100 14.800 ;
        RECT 180.600 14.200 180.900 17.800 ;
        RECT 181.400 15.200 181.700 26.800 ;
        RECT 183.000 26.200 183.300 31.800 ;
        RECT 183.000 25.800 183.400 26.200 ;
        RECT 182.200 22.800 182.600 23.200 ;
        RECT 184.600 23.100 185.000 28.900 ;
        RECT 181.400 14.800 181.800 15.200 ;
        RECT 180.600 13.800 181.000 14.200 ;
        RECT 182.200 13.200 182.500 22.800 ;
        RECT 185.400 17.200 185.700 34.800 ;
        RECT 187.800 32.100 188.200 37.900 ;
        RECT 189.400 35.800 189.800 36.200 ;
        RECT 189.400 35.200 189.700 35.800 ;
        RECT 188.600 34.800 189.000 35.200 ;
        RECT 189.400 34.800 189.800 35.200 ;
        RECT 188.600 34.200 188.900 34.800 ;
        RECT 188.600 33.800 189.000 34.200 ;
        RECT 187.000 29.800 187.400 30.200 ;
        RECT 186.200 25.100 186.600 27.900 ;
        RECT 187.000 26.200 187.300 29.800 ;
        RECT 191.800 29.200 192.100 41.800 ;
        RECT 192.600 32.100 193.000 37.900 ;
        RECT 194.200 37.200 194.500 53.800 ;
        RECT 199.000 52.800 199.400 53.200 ;
        RECT 202.200 53.100 202.600 53.200 ;
        RECT 203.000 53.100 203.400 53.200 ;
        RECT 202.200 52.800 203.400 53.100 ;
        RECT 195.800 51.800 196.200 52.200 ;
        RECT 195.000 47.800 195.400 48.200 ;
        RECT 195.000 39.200 195.300 47.800 ;
        RECT 195.800 46.200 196.100 51.800 ;
        RECT 195.800 45.800 196.200 46.200 ;
        RECT 197.400 43.100 197.800 48.900 ;
        RECT 199.000 47.200 199.300 52.800 ;
        RECT 203.000 52.100 203.400 52.200 ;
        RECT 203.000 51.800 204.100 52.100 ;
        RECT 201.400 49.800 201.800 50.200 ;
        RECT 201.400 49.200 201.700 49.800 ;
        RECT 201.400 48.800 201.800 49.200 ;
        RECT 202.200 48.100 202.600 48.200 ;
        RECT 203.000 48.100 203.400 48.200 ;
        RECT 202.200 47.800 203.400 48.100 ;
        RECT 199.000 46.800 199.400 47.200 ;
        RECT 202.200 47.100 202.600 47.200 ;
        RECT 203.000 47.100 203.400 47.200 ;
        RECT 202.200 46.800 203.400 47.100 ;
        RECT 203.800 46.200 204.100 51.800 ;
        RECT 204.600 46.200 204.900 53.800 ;
        RECT 200.600 45.800 201.000 46.200 ;
        RECT 201.400 45.800 201.800 46.200 ;
        RECT 203.800 45.800 204.200 46.200 ;
        RECT 204.600 45.800 205.000 46.200 ;
        RECT 198.200 43.800 198.600 44.200 ;
        RECT 195.000 38.800 195.400 39.200 ;
        RECT 195.800 38.800 196.200 39.200 ;
        RECT 194.200 36.800 194.600 37.200 ;
        RECT 194.200 33.100 194.600 35.900 ;
        RECT 191.800 28.800 192.200 29.200 ;
        RECT 187.800 27.800 188.200 28.200 ;
        RECT 192.600 28.100 193.000 28.200 ;
        RECT 193.400 28.100 193.800 28.200 ;
        RECT 192.600 27.800 193.800 28.100 ;
        RECT 194.200 28.100 194.600 28.200 ;
        RECT 194.200 27.800 195.300 28.100 ;
        RECT 187.800 26.200 188.100 27.800 ;
        RECT 190.200 26.800 190.600 27.200 ;
        RECT 192.600 26.800 193.000 27.200 ;
        RECT 190.200 26.200 190.500 26.800 ;
        RECT 192.600 26.200 192.900 26.800 ;
        RECT 187.000 25.800 187.400 26.200 ;
        RECT 187.800 25.800 188.200 26.200 ;
        RECT 190.200 25.800 190.600 26.200 ;
        RECT 192.600 25.800 193.000 26.200 ;
        RECT 194.200 25.800 194.600 26.200 ;
        RECT 194.200 25.200 194.500 25.800 ;
        RECT 194.200 24.800 194.600 25.200 ;
        RECT 189.400 21.800 189.800 22.200 ;
        RECT 189.400 19.100 189.700 21.800 ;
        RECT 195.000 19.200 195.300 27.800 ;
        RECT 195.800 26.200 196.100 38.800 ;
        RECT 197.400 32.100 197.800 37.900 ;
        RECT 198.200 35.200 198.500 43.800 ;
        RECT 198.200 34.800 198.600 35.200 ;
        RECT 197.400 30.800 197.800 31.200 ;
        RECT 195.800 25.800 196.200 26.200 ;
        RECT 195.800 22.200 196.100 25.800 ;
        RECT 195.800 21.800 196.200 22.200 ;
        RECT 196.600 21.800 197.000 22.200 ;
        RECT 196.600 20.100 196.900 21.800 ;
        RECT 195.800 19.800 196.900 20.100 ;
        RECT 189.400 18.800 190.500 19.100 ;
        RECT 195.000 18.800 195.400 19.200 ;
        RECT 185.400 16.800 185.800 17.200 ;
        RECT 187.000 16.800 187.400 17.200 ;
        RECT 187.000 15.200 187.300 16.800 ;
        RECT 183.000 15.100 183.400 15.200 ;
        RECT 183.800 15.100 184.200 15.200 ;
        RECT 183.000 14.800 184.200 15.100 ;
        RECT 186.200 14.800 186.600 15.200 ;
        RECT 187.000 14.800 187.400 15.200 ;
        RECT 186.200 14.200 186.500 14.800 ;
        RECT 186.200 13.800 186.600 14.200 ;
        RECT 176.600 12.800 177.000 13.200 ;
        RECT 182.200 13.100 182.600 13.200 ;
        RECT 187.800 13.100 188.200 15.900 ;
        RECT 188.600 13.800 189.000 14.200 ;
        RECT 182.200 12.800 183.300 13.100 ;
        RECT 176.600 11.200 176.900 12.800 ;
        RECT 179.800 11.800 180.200 12.200 ;
        RECT 176.600 10.800 177.000 11.200 ;
        RECT 175.800 9.800 176.900 10.100 ;
        RECT 167.800 6.100 168.200 6.200 ;
        RECT 167.000 5.800 168.200 6.100 ;
        RECT 171.000 3.100 171.400 8.900 ;
        RECT 173.400 8.800 173.800 9.200 ;
        RECT 171.800 7.800 172.200 8.200 ;
        RECT 171.800 7.200 172.100 7.800 ;
        RECT 171.800 6.800 172.200 7.200 ;
        RECT 172.600 5.100 173.000 7.900 ;
        RECT 175.800 3.100 176.200 8.900 ;
        RECT 176.600 7.200 176.900 9.800 ;
        RECT 176.600 6.800 177.000 7.200 ;
        RECT 176.600 6.200 176.900 6.800 ;
        RECT 179.800 6.300 180.100 11.800 ;
        RECT 183.000 9.200 183.300 12.800 ;
        RECT 185.400 12.100 185.800 12.200 ;
        RECT 186.200 12.100 186.600 12.200 ;
        RECT 185.400 11.800 186.600 12.100 ;
        RECT 187.000 11.800 187.400 12.200 ;
        RECT 176.600 5.800 177.000 6.200 ;
        RECT 179.800 5.900 180.200 6.300 ;
        RECT 180.600 3.100 181.000 8.900 ;
        RECT 183.000 8.800 183.400 9.200 ;
        RECT 182.200 5.100 182.600 7.900 ;
        RECT 185.400 3.100 185.800 8.900 ;
        RECT 186.200 6.800 186.600 7.200 ;
        RECT 186.200 6.200 186.500 6.800 ;
        RECT 187.000 6.200 187.300 11.800 ;
        RECT 188.600 7.200 188.900 13.800 ;
        RECT 189.400 12.100 189.800 17.900 ;
        RECT 190.200 15.100 190.500 18.800 ;
        RECT 190.200 14.700 190.600 15.100 ;
        RECT 194.200 12.100 194.600 17.900 ;
        RECT 188.600 6.800 189.000 7.200 ;
        RECT 186.200 5.800 186.600 6.200 ;
        RECT 187.000 5.800 187.400 6.200 ;
        RECT 190.200 3.100 190.600 8.900 ;
        RECT 191.800 5.100 192.200 7.900 ;
        RECT 192.600 5.100 193.000 7.900 ;
        RECT 194.200 3.100 194.600 8.900 ;
        RECT 195.800 6.200 196.100 19.800 ;
        RECT 196.600 18.800 197.000 19.200 ;
        RECT 196.600 18.200 196.900 18.800 ;
        RECT 196.600 17.800 197.000 18.200 ;
        RECT 197.400 15.200 197.700 30.800 ;
        RECT 198.200 26.800 198.600 27.200 ;
        RECT 198.200 26.200 198.500 26.800 ;
        RECT 198.200 25.800 198.600 26.200 ;
        RECT 197.400 14.800 197.800 15.200 ;
        RECT 198.200 9.200 198.500 25.800 ;
        RECT 199.000 21.800 199.400 22.200 ;
        RECT 199.000 19.100 199.300 21.800 ;
        RECT 199.800 19.100 200.200 19.200 ;
        RECT 199.000 18.800 200.200 19.100 ;
        RECT 200.600 15.200 200.900 45.800 ;
        RECT 201.400 35.100 201.700 45.800 ;
        RECT 201.400 34.700 201.800 35.100 ;
        RECT 201.400 32.800 201.800 33.200 ;
        RECT 201.400 26.200 201.700 32.800 ;
        RECT 202.200 32.100 202.600 37.900 ;
        RECT 203.800 33.100 204.200 35.900 ;
        RECT 201.400 25.800 201.800 26.200 ;
        RECT 202.200 26.100 202.600 26.200 ;
        RECT 203.000 26.100 203.400 26.200 ;
        RECT 202.200 25.800 203.400 26.100 ;
        RECT 200.600 14.800 201.000 15.200 ;
        RECT 200.600 12.800 201.000 13.200 ;
        RECT 198.200 8.800 198.600 9.200 ;
        RECT 195.800 5.800 196.200 6.200 ;
        RECT 199.000 3.100 199.400 8.900 ;
        RECT 200.600 7.200 200.900 12.800 ;
        RECT 202.200 9.100 202.600 9.200 ;
        RECT 203.000 9.100 203.400 9.200 ;
        RECT 202.200 8.800 203.400 9.100 ;
        RECT 200.600 6.800 201.000 7.200 ;
      LAYER via2 ;
        RECT 16.600 165.800 17.000 166.200 ;
        RECT 11.800 145.800 12.200 146.200 ;
        RECT 13.400 125.800 13.800 126.200 ;
        RECT 12.600 106.800 13.000 107.200 ;
        RECT 27.800 124.800 28.200 125.200 ;
        RECT 20.600 114.800 21.000 115.200 ;
        RECT 24.600 106.800 25.000 107.200 ;
        RECT 13.400 105.800 13.800 106.200 ;
        RECT 12.600 94.800 13.000 95.200 ;
        RECT 23.000 95.800 23.400 96.200 ;
        RECT 19.800 94.800 20.200 95.200 ;
        RECT 5.400 74.800 5.800 75.200 ;
        RECT 13.400 74.800 13.800 75.200 ;
        RECT 16.600 74.800 17.000 75.200 ;
        RECT 5.400 65.800 5.800 66.200 ;
        RECT 1.400 34.800 1.800 35.200 ;
        RECT 10.200 68.800 10.600 69.200 ;
        RECT 14.200 66.800 14.600 67.200 ;
        RECT 11.800 65.800 12.200 66.200 ;
        RECT 11.800 38.800 12.200 39.200 ;
        RECT 51.800 165.800 52.200 166.200 ;
        RECT 36.600 125.800 37.000 126.200 ;
        RECT 52.600 154.800 53.000 155.200 ;
        RECT 57.400 155.800 57.800 156.200 ;
        RECT 54.200 147.800 54.600 148.200 ;
        RECT 59.000 153.800 59.400 154.200 ;
        RECT 67.800 165.800 68.200 166.200 ;
        RECT 42.200 134.800 42.600 135.200 ;
        RECT 30.200 114.800 30.600 115.200 ;
        RECT 56.600 134.800 57.000 135.200 ;
        RECT 47.800 126.800 48.200 127.200 ;
        RECT 42.200 113.800 42.600 114.200 ;
        RECT 59.800 127.800 60.200 128.200 ;
        RECT 59.000 126.800 59.400 127.200 ;
        RECT 85.400 173.800 85.800 174.200 ;
        RECT 74.200 155.800 74.600 156.200 ;
        RECT 77.400 153.800 77.800 154.200 ;
        RECT 97.400 168.800 97.800 169.200 ;
        RECT 123.000 172.800 123.400 173.200 ;
        RECT 104.600 166.800 105.000 167.200 ;
        RECT 89.400 146.800 89.800 147.200 ;
        RECT 67.000 126.800 67.400 127.200 ;
        RECT 48.600 113.800 49.000 114.200 ;
        RECT 31.800 107.800 32.200 108.200 ;
        RECT 30.200 106.800 30.600 107.200 ;
        RECT 35.000 106.800 35.400 107.200 ;
        RECT 27.000 105.800 27.400 106.200 ;
        RECT 32.600 105.800 33.000 106.200 ;
        RECT 40.600 107.800 41.000 108.200 ;
        RECT 46.200 107.800 46.600 108.200 ;
        RECT 60.600 113.800 61.000 114.200 ;
        RECT 63.800 113.800 64.200 114.200 ;
        RECT 37.400 106.800 37.800 107.200 ;
        RECT 42.200 106.800 42.600 107.200 ;
        RECT 51.800 105.800 52.200 106.200 ;
        RECT 27.000 92.800 27.400 93.200 ;
        RECT 39.000 86.800 39.400 87.200 ;
        RECT 26.200 66.800 26.600 67.200 ;
        RECT 36.600 74.800 37.000 75.200 ;
        RECT 30.200 65.800 30.600 66.200 ;
        RECT 32.600 65.800 33.000 66.200 ;
        RECT 21.400 56.800 21.800 57.200 ;
        RECT 23.000 44.800 23.400 45.200 ;
        RECT 17.400 33.800 17.800 34.200 ;
        RECT 14.200 14.800 14.600 15.200 ;
        RECT 27.800 45.900 28.200 46.300 ;
        RECT 32.600 64.800 33.000 65.200 ;
        RECT 30.200 54.800 30.600 55.200 ;
        RECT 37.400 65.800 37.800 66.200 ;
        RECT 48.600 93.800 49.000 94.200 ;
        RECT 50.200 88.800 50.600 89.200 ;
        RECT 59.000 93.800 59.400 94.200 ;
        RECT 124.600 167.800 125.000 168.200 ;
        RECT 107.000 154.800 107.400 155.200 ;
        RECT 117.400 163.800 117.800 164.200 ;
        RECT 112.600 154.800 113.000 155.200 ;
        RECT 115.000 144.800 115.400 145.200 ;
        RECT 90.200 128.800 90.600 129.200 ;
        RECT 88.600 127.800 89.000 128.200 ;
        RECT 83.000 124.800 83.400 125.200 ;
        RECT 86.200 125.800 86.600 126.200 ;
        RECT 69.400 105.800 69.800 106.200 ;
        RECT 66.200 94.800 66.600 95.200 ;
        RECT 64.600 93.800 65.000 94.200 ;
        RECT 79.000 94.800 79.400 95.200 ;
        RECT 85.400 108.800 85.800 109.200 ;
        RECT 97.400 133.800 97.800 134.200 ;
        RECT 90.200 107.800 90.600 108.200 ;
        RECT 93.400 106.800 93.800 107.200 ;
        RECT 96.600 105.800 97.000 106.200 ;
        RECT 91.000 104.800 91.400 105.200 ;
        RECT 85.400 94.800 85.800 95.200 ;
        RECT 61.400 84.800 61.800 85.200 ;
        RECT 44.600 75.800 45.000 76.200 ;
        RECT 51.000 75.800 51.400 76.200 ;
        RECT 47.000 74.800 47.400 75.200 ;
        RECT 50.200 67.800 50.600 68.200 ;
        RECT 52.600 66.800 53.000 67.200 ;
        RECT 42.200 63.800 42.600 64.200 ;
        RECT 37.400 55.800 37.800 56.200 ;
        RECT 27.800 34.800 28.200 35.200 ;
        RECT 37.400 46.800 37.800 47.200 ;
        RECT 35.000 34.800 35.400 35.200 ;
        RECT 19.800 14.800 20.200 15.200 ;
        RECT 74.200 85.800 74.600 86.200 ;
        RECT 77.400 85.800 77.800 86.200 ;
        RECT 71.800 84.800 72.200 85.200 ;
        RECT 83.800 92.800 84.200 93.200 ;
        RECT 73.400 74.800 73.800 75.200 ;
        RECT 79.000 74.800 79.400 75.200 ;
        RECT 66.200 73.800 66.600 74.200 ;
        RECT 59.000 68.800 59.400 69.200 ;
        RECT 55.800 64.800 56.200 65.200 ;
        RECT 56.600 56.800 57.000 57.200 ;
        RECT 46.200 35.800 46.600 36.200 ;
        RECT 32.600 27.800 33.000 28.200 ;
        RECT 25.400 16.800 25.800 17.200 ;
        RECT 29.400 15.800 29.800 16.200 ;
        RECT 27.800 14.800 28.200 15.200 ;
        RECT 38.200 18.800 38.600 19.200 ;
        RECT 45.400 26.800 45.800 27.200 ;
        RECT 46.200 25.800 46.600 26.200 ;
        RECT 48.600 24.800 49.000 25.200 ;
        RECT 26.200 13.800 26.600 14.200 ;
        RECT 31.800 13.800 32.200 14.200 ;
        RECT 19.000 5.800 19.400 6.200 ;
        RECT 44.600 14.800 45.000 15.200 ;
        RECT 50.200 17.800 50.600 18.200 ;
        RECT 68.600 72.800 69.000 73.200 ;
        RECT 70.200 67.800 70.600 68.200 ;
        RECT 71.000 65.800 71.400 66.200 ;
        RECT 63.800 53.800 64.200 54.200 ;
        RECT 71.000 54.800 71.400 55.200 ;
        RECT 59.800 35.800 60.200 36.200 ;
        RECT 76.600 57.800 77.000 58.200 ;
        RECT 63.800 35.800 64.200 36.200 ;
        RECT 66.200 33.800 66.600 34.200 ;
        RECT 93.400 94.800 93.800 95.200 ;
        RECT 90.200 88.800 90.600 89.200 ;
        RECT 87.800 86.800 88.200 87.200 ;
        RECT 92.600 86.800 93.000 87.200 ;
        RECT 84.600 66.800 85.000 67.200 ;
        RECT 88.600 71.800 89.000 72.200 ;
        RECT 93.400 74.800 93.800 75.200 ;
        RECT 109.400 134.800 109.800 135.200 ;
        RECT 105.400 125.800 105.800 126.200 ;
        RECT 122.200 145.800 122.600 146.200 ;
        RECT 123.000 143.800 123.400 144.200 ;
        RECT 132.600 163.800 133.000 164.200 ;
        RECT 143.800 151.800 144.200 152.200 ;
        RECT 131.000 147.800 131.400 148.200 ;
        RECT 137.400 146.800 137.800 147.200 ;
        RECT 126.200 143.800 126.600 144.200 ;
        RECT 107.800 131.800 108.200 132.200 ;
        RECT 107.800 126.800 108.200 127.200 ;
        RECT 117.400 122.800 117.800 123.200 ;
        RECT 105.400 113.800 105.800 114.200 ;
        RECT 118.200 113.800 118.600 114.200 ;
        RECT 193.400 172.800 193.800 173.200 ;
        RECT 201.400 172.800 201.800 173.200 ;
        RECT 183.800 166.800 184.200 167.200 ;
        RECT 151.800 147.800 152.200 148.200 ;
        RECT 161.400 147.800 161.800 148.200 ;
        RECT 131.000 134.800 131.400 135.200 ;
        RECT 138.200 134.800 138.600 135.200 ;
        RECT 96.600 74.800 97.000 75.200 ;
        RECT 93.400 66.800 93.800 67.200 ;
        RECT 99.000 66.800 99.400 67.200 ;
        RECT 96.600 64.800 97.000 65.200 ;
        RECT 55.000 25.800 55.400 26.200 ;
        RECT 61.400 29.800 61.800 30.200 ;
        RECT 73.400 25.800 73.800 26.200 ;
        RECT 72.600 24.800 73.000 25.200 ;
        RECT 47.000 5.800 47.400 6.200 ;
        RECT 58.200 5.800 58.600 6.200 ;
        RECT 95.000 48.800 95.400 49.200 ;
        RECT 117.400 102.800 117.800 103.200 ;
        RECT 115.800 94.800 116.200 95.200 ;
        RECT 72.600 13.800 73.000 14.200 ;
        RECT 79.800 14.800 80.200 15.200 ;
        RECT 66.200 4.800 66.600 5.200 ;
        RECT 87.000 33.800 87.400 34.200 ;
        RECT 130.200 114.800 130.600 115.200 ;
        RECT 119.800 95.800 120.200 96.200 ;
        RECT 131.800 108.800 132.200 109.200 ;
        RECT 132.600 106.800 133.000 107.200 ;
        RECT 123.000 93.800 123.400 94.200 ;
        RECT 119.000 85.800 119.400 86.200 ;
        RECT 115.000 78.800 115.400 79.200 ;
        RECT 116.600 74.800 117.000 75.200 ;
        RECT 119.800 76.800 120.200 77.200 ;
        RECT 137.400 128.800 137.800 129.200 ;
        RECT 138.200 126.800 138.600 127.200 ;
        RECT 147.000 144.800 147.400 145.200 ;
        RECT 149.400 135.800 149.800 136.200 ;
        RECT 170.200 148.800 170.600 149.200 ;
        RECT 164.600 134.800 165.000 135.200 ;
        RECT 145.400 128.800 145.800 129.200 ;
        RECT 139.000 125.800 139.400 126.200 ;
        RECT 137.400 105.800 137.800 106.200 ;
        RECT 131.800 86.800 132.200 87.200 ;
        RECT 162.200 127.800 162.600 128.200 ;
        RECT 162.200 126.800 162.600 127.200 ;
        RECT 158.200 125.800 158.600 126.200 ;
        RECT 179.000 135.800 179.400 136.200 ;
        RECT 187.000 145.800 187.400 146.200 ;
        RECT 187.000 143.800 187.400 144.200 ;
        RECT 183.800 134.800 184.200 135.200 ;
        RECT 169.400 126.800 169.800 127.200 ;
        RECT 167.800 125.800 168.200 126.200 ;
        RECT 165.400 124.800 165.800 125.200 ;
        RECT 192.600 133.800 193.000 134.200 ;
        RECT 196.600 133.800 197.000 134.200 ;
        RECT 203.000 127.800 203.400 128.200 ;
        RECT 187.800 126.800 188.200 127.200 ;
        RECT 194.200 125.800 194.600 126.200 ;
        RECT 171.800 124.800 172.200 125.200 ;
        RECT 164.600 115.800 165.000 116.200 ;
        RECT 157.400 113.800 157.800 114.200 ;
        RECT 111.000 65.800 111.400 66.200 ;
        RECT 119.800 67.800 120.200 68.200 ;
        RECT 116.600 54.800 117.000 55.200 ;
        RECT 107.800 46.800 108.200 47.200 ;
        RECT 112.600 46.800 113.000 47.200 ;
        RECT 135.000 72.800 135.400 73.200 ;
        RECT 107.000 45.800 107.400 46.200 ;
        RECT 112.600 45.800 113.000 46.200 ;
        RECT 94.200 26.800 94.600 27.200 ;
        RECT 93.400 25.800 93.800 26.200 ;
        RECT 86.200 15.800 86.600 16.200 ;
        RECT 82.200 13.800 82.600 14.200 ;
        RECT 113.400 44.800 113.800 45.200 ;
        RECT 109.400 36.800 109.800 37.200 ;
        RECT 113.400 33.800 113.800 34.200 ;
        RECT 152.600 93.800 153.000 94.200 ;
        RECT 151.000 92.800 151.400 93.200 ;
        RECT 155.000 92.800 155.400 93.200 ;
        RECT 159.800 92.800 160.200 93.200 ;
        RECT 173.400 108.800 173.800 109.200 ;
        RECT 169.400 107.800 169.800 108.200 ;
        RECT 176.600 107.800 177.000 108.200 ;
        RECT 149.400 85.800 149.800 86.200 ;
        RECT 151.800 85.800 152.200 86.200 ;
        RECT 147.800 84.800 148.200 85.200 ;
        RECT 139.800 72.800 140.200 73.200 ;
        RECT 131.000 65.800 131.400 66.200 ;
        RECT 129.400 53.800 129.800 54.200 ;
        RECT 103.000 8.800 103.400 9.200 ;
        RECT 135.000 48.800 135.400 49.200 ;
        RECT 145.400 67.800 145.800 68.200 ;
        RECT 155.000 73.800 155.400 74.200 ;
        RECT 158.200 73.800 158.600 74.200 ;
        RECT 147.800 64.800 148.200 65.200 ;
        RECT 142.200 53.800 142.600 54.200 ;
        RECT 151.000 54.800 151.400 55.200 ;
        RECT 128.600 34.800 129.000 35.200 ;
        RECT 125.400 26.800 125.800 27.200 ;
        RECT 130.200 31.800 130.600 32.200 ;
        RECT 150.200 47.800 150.600 48.200 ;
        RECT 127.800 26.800 128.200 27.200 ;
        RECT 133.400 26.800 133.800 27.200 ;
        RECT 120.600 25.800 121.000 26.200 ;
        RECT 124.600 25.800 125.000 26.200 ;
        RECT 127.000 25.800 127.400 26.200 ;
        RECT 120.600 24.800 121.000 25.200 ;
        RECT 119.000 14.800 119.400 15.200 ;
        RECT 133.400 8.800 133.800 9.200 ;
        RECT 144.600 25.800 145.000 26.200 ;
        RECT 180.600 95.800 181.000 96.200 ;
        RECT 197.400 106.800 197.800 107.200 ;
        RECT 191.000 105.800 191.400 106.200 ;
        RECT 177.400 85.800 177.800 86.200 ;
        RECT 179.000 73.800 179.400 74.200 ;
        RECT 165.400 63.800 165.800 64.200 ;
        RECT 168.600 64.800 169.000 65.200 ;
        RECT 195.000 104.800 195.400 105.200 ;
        RECT 195.000 85.800 195.400 86.200 ;
        RECT 195.800 74.800 196.200 75.200 ;
        RECT 194.200 73.800 194.600 74.200 ;
        RECT 174.200 41.800 174.600 42.200 ;
        RECT 192.600 55.800 193.000 56.200 ;
        RECT 188.600 47.800 189.000 48.200 ;
        RECT 195.800 72.800 196.200 73.200 ;
        RECT 200.600 55.800 201.000 56.200 ;
        RECT 187.800 45.800 188.200 46.200 ;
        RECT 159.800 27.800 160.200 28.200 ;
        RECT 164.600 25.800 165.000 26.200 ;
        RECT 146.200 13.800 146.600 14.200 ;
        RECT 153.400 8.800 153.800 9.200 ;
        RECT 203.000 52.800 203.400 53.200 ;
        RECT 203.000 46.800 203.400 47.200 ;
        RECT 186.200 11.800 186.600 12.200 ;
        RECT 203.000 25.800 203.400 26.200 ;
      LAYER metal3 ;
        RECT 196.600 177.100 197.000 177.200 ;
        RECT 195.000 176.800 197.000 177.100 ;
        RECT 195.000 176.200 195.300 176.800 ;
        RECT 195.000 175.800 195.400 176.200 ;
        RECT 60.600 175.100 61.000 175.200 ;
        RECT 67.000 175.100 67.400 175.200 ;
        RECT 60.600 174.800 67.400 175.100 ;
        RECT 79.800 174.800 80.200 175.200 ;
        RECT 35.000 174.100 35.400 174.200 ;
        RECT 37.400 174.100 37.800 174.200 ;
        RECT 35.000 173.800 37.800 174.100 ;
        RECT 65.400 174.100 65.800 174.200 ;
        RECT 77.400 174.100 77.800 174.200 ;
        RECT 65.400 173.800 77.800 174.100 ;
        RECT 79.800 174.100 80.100 174.800 ;
        RECT 85.400 174.100 85.800 174.200 ;
        RECT 79.800 173.800 85.800 174.100 ;
        RECT 91.000 174.100 91.400 174.200 ;
        RECT 94.200 174.100 94.600 174.200 ;
        RECT 91.000 173.800 94.600 174.100 ;
        RECT 100.600 173.800 101.000 174.200 ;
        RECT 114.200 174.100 114.600 174.200 ;
        RECT 135.000 174.100 135.400 174.200 ;
        RECT 114.200 173.800 135.400 174.100 ;
        RECT 139.000 173.800 139.400 174.200 ;
        RECT 146.200 174.100 146.600 174.200 ;
        RECT 148.600 174.100 149.000 174.200 ;
        RECT 151.000 174.100 151.400 174.200 ;
        RECT 146.200 173.800 151.400 174.100 ;
        RECT 157.400 173.800 157.800 174.200 ;
        RECT 182.200 173.800 182.600 174.200 ;
        RECT 195.000 173.800 195.400 174.200 ;
        RECT 66.200 173.100 66.600 173.200 ;
        RECT 53.400 172.800 66.600 173.100 ;
        RECT 92.600 173.100 93.000 173.200 ;
        RECT 100.600 173.100 100.900 173.800 ;
        RECT 115.000 173.100 115.400 173.200 ;
        RECT 92.600 172.800 115.400 173.100 ;
        RECT 121.400 173.100 121.800 173.200 ;
        RECT 123.000 173.100 123.400 173.200 ;
        RECT 129.400 173.100 129.800 173.200 ;
        RECT 121.400 172.800 129.800 173.100 ;
        RECT 139.000 173.100 139.300 173.800 ;
        RECT 143.800 173.100 144.200 173.200 ;
        RECT 151.000 173.100 151.400 173.200 ;
        RECT 157.400 173.100 157.700 173.800 ;
        RECT 173.400 173.100 173.800 173.200 ;
        RECT 182.200 173.100 182.500 173.800 ;
        RECT 139.000 172.800 182.500 173.100 ;
        RECT 193.400 173.100 193.800 173.200 ;
        RECT 195.000 173.100 195.300 173.800 ;
        RECT 193.400 172.800 195.300 173.100 ;
        RECT 196.600 172.800 197.000 173.200 ;
        RECT 201.400 173.100 201.800 173.200 ;
        RECT 202.200 173.100 202.600 173.200 ;
        RECT 201.400 172.800 202.600 173.100 ;
        RECT 53.400 172.200 53.700 172.800 ;
        RECT 196.600 172.200 196.900 172.800 ;
        RECT 44.600 172.100 45.000 172.200 ;
        RECT 53.400 172.100 53.800 172.200 ;
        RECT 44.600 171.800 53.800 172.100 ;
        RECT 68.600 172.100 69.000 172.200 ;
        RECT 71.000 172.100 71.400 172.200 ;
        RECT 68.600 171.800 71.400 172.100 ;
        RECT 82.200 172.100 82.600 172.200 ;
        RECT 111.800 172.100 112.200 172.200 ;
        RECT 82.200 171.800 112.200 172.100 ;
        RECT 119.000 172.100 119.400 172.200 ;
        RECT 122.200 172.100 122.600 172.200 ;
        RECT 119.000 171.800 122.600 172.100 ;
        RECT 190.200 171.800 190.600 172.200 ;
        RECT 196.600 171.800 197.000 172.200 ;
        RECT 190.200 171.200 190.500 171.800 ;
        RECT 49.400 171.100 49.800 171.200 ;
        RECT 51.000 171.100 51.400 171.200 ;
        RECT 49.400 170.800 51.400 171.100 ;
        RECT 57.400 171.100 57.800 171.200 ;
        RECT 82.200 171.100 82.600 171.200 ;
        RECT 57.400 170.800 82.600 171.100 ;
        RECT 190.200 170.800 190.600 171.200 ;
        RECT 14.200 170.100 14.600 170.200 ;
        RECT 19.000 170.100 19.400 170.200 ;
        RECT 14.200 169.800 19.400 170.100 ;
        RECT 30.200 170.100 30.600 170.200 ;
        RECT 48.600 170.100 49.000 170.200 ;
        RECT 30.200 169.800 49.000 170.100 ;
        RECT 126.200 170.100 126.600 170.200 ;
        RECT 140.600 170.100 141.000 170.200 ;
        RECT 126.200 169.800 141.000 170.100 ;
        RECT 9.400 168.800 9.800 169.200 ;
        RECT 16.600 169.100 17.000 169.200 ;
        RECT 35.800 169.100 36.200 169.200 ;
        RECT 16.600 168.800 36.200 169.100 ;
        RECT 97.400 169.100 97.800 169.200 ;
        RECT 99.000 169.100 99.400 169.200 ;
        RECT 97.400 168.800 99.400 169.100 ;
        RECT 161.400 169.100 161.800 169.200 ;
        RECT 167.000 169.100 167.400 169.200 ;
        RECT 161.400 168.800 167.400 169.100 ;
        RECT 180.600 169.100 181.000 169.200 ;
        RECT 184.600 169.100 185.000 169.200 ;
        RECT 180.600 168.800 185.000 169.100 ;
        RECT 190.200 168.800 190.600 169.200 ;
        RECT 203.800 168.800 204.200 169.200 ;
        RECT 9.400 168.100 9.700 168.800 ;
        RECT 11.000 168.100 11.400 168.200 ;
        RECT 28.600 168.100 29.000 168.200 ;
        RECT 9.400 167.800 29.000 168.100 ;
        RECT 99.000 168.100 99.400 168.200 ;
        RECT 100.600 168.100 101.000 168.200 ;
        RECT 106.200 168.100 106.600 168.200 ;
        RECT 109.400 168.100 109.800 168.200 ;
        RECT 99.000 167.800 109.800 168.100 ;
        RECT 124.600 168.100 125.000 168.200 ;
        RECT 125.400 168.100 125.800 168.200 ;
        RECT 134.200 168.100 134.600 168.200 ;
        RECT 124.600 167.800 134.600 168.100 ;
        RECT 187.800 168.100 188.200 168.200 ;
        RECT 190.200 168.100 190.500 168.800 ;
        RECT 187.800 167.800 190.500 168.100 ;
        RECT 198.200 168.100 198.600 168.200 ;
        RECT 203.800 168.100 204.100 168.800 ;
        RECT 198.200 167.800 204.100 168.100 ;
        RECT 39.800 167.100 40.200 167.200 ;
        RECT 57.400 167.100 57.800 167.200 ;
        RECT 39.800 166.800 57.800 167.100 ;
        RECT 81.400 167.100 81.800 167.200 ;
        RECT 90.200 167.100 90.600 167.200 ;
        RECT 81.400 166.800 90.600 167.100 ;
        RECT 104.600 167.100 105.000 167.200 ;
        RECT 107.000 167.100 107.400 167.200 ;
        RECT 104.600 166.800 107.400 167.100 ;
        RECT 115.800 167.100 116.200 167.200 ;
        RECT 117.400 167.100 117.800 167.200 ;
        RECT 124.600 167.100 125.000 167.200 ;
        RECT 115.800 166.800 125.000 167.100 ;
        RECT 125.400 167.100 125.800 167.200 ;
        RECT 128.600 167.100 129.000 167.200 ;
        RECT 155.000 167.100 155.400 167.200 ;
        RECT 125.400 166.800 129.000 167.100 ;
        RECT 154.200 166.800 155.400 167.100 ;
        RECT 183.800 167.100 184.200 167.200 ;
        RECT 190.200 167.100 190.600 167.200 ;
        RECT 191.000 167.100 191.400 167.200 ;
        RECT 204.600 167.100 205.000 167.200 ;
        RECT 183.800 166.800 205.000 167.100 ;
        RECT 154.200 166.200 154.500 166.800 ;
        RECT 16.600 166.100 17.000 166.200 ;
        RECT 23.000 166.100 23.400 166.200 ;
        RECT 16.600 165.800 23.400 166.100 ;
        RECT 51.800 166.100 52.200 166.200 ;
        RECT 53.400 166.100 53.800 166.200 ;
        RECT 51.800 165.800 53.800 166.100 ;
        RECT 64.600 166.100 65.000 166.200 ;
        RECT 67.800 166.100 68.200 166.200 ;
        RECT 111.000 166.100 111.400 166.200 ;
        RECT 112.600 166.100 113.000 166.200 ;
        RECT 64.600 165.800 113.000 166.100 ;
        RECT 114.200 166.100 114.600 166.200 ;
        RECT 118.200 166.100 118.600 166.200 ;
        RECT 114.200 165.800 118.600 166.100 ;
        RECT 120.600 166.100 121.000 166.200 ;
        RECT 128.600 166.100 129.000 166.200 ;
        RECT 120.600 165.800 129.000 166.100 ;
        RECT 154.200 165.800 154.600 166.200 ;
        RECT 159.000 166.100 159.400 166.200 ;
        RECT 161.400 166.100 161.800 166.200 ;
        RECT 159.000 165.800 161.800 166.100 ;
        RECT 189.400 166.100 189.800 166.200 ;
        RECT 199.000 166.100 199.400 166.200 ;
        RECT 189.400 165.800 199.400 166.100 ;
        RECT 201.400 165.800 201.800 166.200 ;
        RECT 201.400 165.200 201.700 165.800 ;
        RECT 35.000 165.100 35.400 165.200 ;
        RECT 58.200 165.100 58.600 165.200 ;
        RECT 66.200 165.100 66.600 165.200 ;
        RECT 79.000 165.100 79.400 165.200 ;
        RECT 35.000 164.800 79.400 165.100 ;
        RECT 94.200 165.100 94.600 165.200 ;
        RECT 111.800 165.100 112.200 165.200 ;
        RECT 94.200 164.800 106.500 165.100 ;
        RECT 98.200 164.200 98.500 164.800 ;
        RECT 106.200 164.200 106.500 164.800 ;
        RECT 108.600 164.800 112.200 165.100 ;
        RECT 121.400 165.100 121.800 165.200 ;
        RECT 125.400 165.100 125.800 165.200 ;
        RECT 121.400 164.800 125.800 165.100 ;
        RECT 179.800 165.100 180.200 165.200 ;
        RECT 183.800 165.100 184.200 165.200 ;
        RECT 187.000 165.100 187.400 165.200 ;
        RECT 179.800 164.800 187.400 165.100 ;
        RECT 197.400 165.100 197.800 165.200 ;
        RECT 199.800 165.100 200.200 165.200 ;
        RECT 197.400 164.800 200.200 165.100 ;
        RECT 201.400 164.800 201.800 165.200 ;
        RECT 108.600 164.200 108.900 164.800 ;
        RECT 28.600 164.100 29.000 164.200 ;
        RECT 71.800 164.100 72.200 164.200 ;
        RECT 28.600 163.800 72.200 164.100 ;
        RECT 98.200 163.800 98.600 164.200 ;
        RECT 106.200 163.800 106.600 164.200 ;
        RECT 108.600 163.800 109.000 164.200 ;
        RECT 117.400 164.100 117.800 164.200 ;
        RECT 120.600 164.100 121.000 164.200 ;
        RECT 117.400 163.800 121.000 164.100 ;
        RECT 132.600 164.100 133.000 164.200 ;
        RECT 145.400 164.100 145.800 164.200 ;
        RECT 132.600 163.800 145.800 164.100 ;
        RECT 164.600 164.100 165.000 164.200 ;
        RECT 165.400 164.100 165.800 164.200 ;
        RECT 196.600 164.100 197.000 164.200 ;
        RECT 197.400 164.100 197.800 164.200 ;
        RECT 164.600 163.800 197.800 164.100 ;
        RECT 46.200 163.100 46.600 163.200 ;
        RECT 73.400 163.100 73.800 163.200 ;
        RECT 46.200 162.800 73.800 163.100 ;
        RECT 107.000 163.100 107.400 163.200 ;
        RECT 116.600 163.100 117.000 163.200 ;
        RECT 107.000 162.800 117.000 163.100 ;
        RECT 24.600 162.100 25.000 162.200 ;
        RECT 59.000 162.100 59.400 162.200 ;
        RECT 61.400 162.100 61.800 162.200 ;
        RECT 71.000 162.100 71.400 162.200 ;
        RECT 24.600 161.800 71.400 162.100 ;
        RECT 75.800 162.100 76.200 162.200 ;
        RECT 79.800 162.100 80.200 162.200 ;
        RECT 82.200 162.100 82.600 162.200 ;
        RECT 115.000 162.100 115.400 162.200 ;
        RECT 75.800 161.800 82.600 162.100 ;
        RECT 103.000 161.800 115.400 162.100 ;
        RECT 123.000 161.800 123.400 162.200 ;
        RECT 103.000 161.200 103.300 161.800 ;
        RECT 123.000 161.200 123.300 161.800 ;
        RECT 75.000 161.100 75.400 161.200 ;
        RECT 78.200 161.100 78.600 161.200 ;
        RECT 75.000 160.800 78.600 161.100 ;
        RECT 103.000 160.800 103.400 161.200 ;
        RECT 123.000 160.800 123.400 161.200 ;
        RECT 55.000 160.100 55.400 160.200 ;
        RECT 77.400 160.100 77.800 160.200 ;
        RECT 55.000 159.800 77.800 160.100 ;
        RECT 169.400 160.100 169.800 160.200 ;
        RECT 171.800 160.100 172.200 160.200 ;
        RECT 169.400 159.800 172.200 160.100 ;
        RECT 63.000 158.800 63.400 159.200 ;
        RECT 83.800 159.100 84.200 159.200 ;
        RECT 84.600 159.100 85.000 159.200 ;
        RECT 83.800 158.800 85.000 159.100 ;
        RECT 121.400 159.100 121.800 159.200 ;
        RECT 124.600 159.100 125.000 159.200 ;
        RECT 121.400 158.800 125.000 159.100 ;
        RECT 63.000 158.200 63.300 158.800 ;
        RECT 63.000 157.800 63.400 158.200 ;
        RECT 97.400 157.800 97.800 158.200 ;
        RECT 112.600 158.100 113.000 158.200 ;
        RECT 116.600 158.100 117.000 158.200 ;
        RECT 127.800 158.100 128.200 158.200 ;
        RECT 112.600 157.800 128.200 158.100 ;
        RECT 173.400 158.100 173.800 158.200 ;
        RECT 195.800 158.100 196.200 158.200 ;
        RECT 173.400 157.800 196.200 158.100 ;
        RECT 52.600 156.800 53.000 157.200 ;
        RECT 75.800 157.100 76.200 157.200 ;
        RECT 61.400 156.800 76.200 157.100 ;
        RECT 77.400 157.100 77.800 157.200 ;
        RECT 97.400 157.100 97.700 157.800 ;
        RECT 77.400 156.800 97.700 157.100 ;
        RECT 108.600 157.100 109.000 157.200 ;
        RECT 114.200 157.100 114.600 157.200 ;
        RECT 108.600 156.800 114.600 157.100 ;
        RECT 115.000 157.100 115.400 157.200 ;
        RECT 117.400 157.100 117.800 157.200 ;
        RECT 115.000 156.800 117.800 157.100 ;
        RECT 184.600 156.800 185.000 157.200 ;
        RECT 4.600 156.100 5.000 156.200 ;
        RECT 21.400 156.100 21.800 156.200 ;
        RECT 4.600 155.800 21.800 156.100 ;
        RECT 43.800 156.100 44.200 156.200 ;
        RECT 52.600 156.100 52.900 156.800 ;
        RECT 61.400 156.200 61.700 156.800 ;
        RECT 43.800 155.800 52.900 156.100 ;
        RECT 57.400 156.100 57.800 156.200 ;
        RECT 61.400 156.100 61.800 156.200 ;
        RECT 57.400 155.800 61.800 156.100 ;
        RECT 63.000 155.800 63.400 156.200 ;
        RECT 71.000 156.100 71.400 156.200 ;
        RECT 74.200 156.100 74.600 156.200 ;
        RECT 115.800 156.100 116.200 156.200 ;
        RECT 71.000 155.800 116.200 156.100 ;
        RECT 119.000 156.100 119.400 156.200 ;
        RECT 129.400 156.100 129.800 156.200 ;
        RECT 119.000 155.800 129.800 156.100 ;
        RECT 179.000 156.100 179.400 156.200 ;
        RECT 184.600 156.100 184.900 156.800 ;
        RECT 179.000 155.800 184.900 156.100 ;
        RECT 190.200 155.800 190.600 156.200 ;
        RECT 3.800 155.100 4.200 155.200 ;
        RECT 17.400 155.100 17.800 155.200 ;
        RECT 3.800 154.800 17.800 155.100 ;
        RECT 21.400 155.100 21.800 155.200 ;
        RECT 52.600 155.100 53.000 155.200 ;
        RECT 56.600 155.100 57.000 155.200 ;
        RECT 21.400 154.800 57.000 155.100 ;
        RECT 59.800 155.100 60.200 155.200 ;
        RECT 63.000 155.100 63.300 155.800 ;
        RECT 59.800 154.800 63.300 155.100 ;
        RECT 84.600 154.800 85.000 155.200 ;
        RECT 106.200 155.100 106.600 155.200 ;
        RECT 107.000 155.100 107.400 155.200 ;
        RECT 106.200 154.800 107.400 155.100 ;
        RECT 111.800 155.100 112.200 155.200 ;
        RECT 112.600 155.100 113.000 155.200 ;
        RECT 111.800 154.800 113.000 155.100 ;
        RECT 158.200 155.100 158.600 155.200 ;
        RECT 162.200 155.100 162.600 155.200 ;
        RECT 158.200 154.800 162.600 155.100 ;
        RECT 180.600 155.100 181.000 155.200 ;
        RECT 188.600 155.100 189.000 155.200 ;
        RECT 190.200 155.100 190.500 155.800 ;
        RECT 180.600 154.800 190.500 155.100 ;
        RECT 44.600 154.100 45.000 154.200 ;
        RECT 59.000 154.100 59.400 154.200 ;
        RECT 64.600 154.100 65.000 154.200 ;
        RECT 44.600 153.800 65.000 154.100 ;
        RECT 77.400 154.100 77.800 154.200 ;
        RECT 84.600 154.100 84.900 154.800 ;
        RECT 77.400 153.800 84.900 154.100 ;
        RECT 95.800 154.100 96.200 154.200 ;
        RECT 100.600 154.100 101.000 154.200 ;
        RECT 104.600 154.100 105.000 154.200 ;
        RECT 95.800 153.800 105.000 154.100 ;
        RECT 110.200 153.800 110.600 154.200 ;
        RECT 113.400 153.800 113.800 154.200 ;
        RECT 115.000 154.100 115.400 154.200 ;
        RECT 121.400 154.100 121.800 154.200 ;
        RECT 115.000 153.800 121.800 154.100 ;
        RECT 133.400 154.100 133.800 154.200 ;
        RECT 151.000 154.100 151.400 154.200 ;
        RECT 151.800 154.100 152.200 154.200 ;
        RECT 133.400 153.800 152.200 154.100 ;
        RECT 169.400 153.800 169.800 154.200 ;
        RECT 183.000 154.100 183.400 154.200 ;
        RECT 188.600 154.100 189.000 154.200 ;
        RECT 183.000 153.800 189.000 154.100 ;
        RECT 189.400 154.100 189.800 154.200 ;
        RECT 190.200 154.100 190.600 154.200 ;
        RECT 189.400 153.800 190.600 154.100 ;
        RECT 13.400 153.100 13.800 153.200 ;
        RECT 14.200 153.100 14.600 153.200 ;
        RECT 16.600 153.100 17.000 153.200 ;
        RECT 35.800 153.100 36.200 153.200 ;
        RECT 38.200 153.100 38.600 153.200 ;
        RECT 110.200 153.100 110.500 153.800 ;
        RECT 13.400 152.800 110.500 153.100 ;
        RECT 113.400 153.100 113.700 153.800 ;
        RECT 138.200 153.100 138.600 153.200 ;
        RECT 147.000 153.100 147.400 153.200 ;
        RECT 113.400 152.800 147.400 153.100 ;
        RECT 169.400 153.100 169.700 153.800 ;
        RECT 173.400 153.100 173.800 153.200 ;
        RECT 175.000 153.100 175.400 153.200 ;
        RECT 169.400 152.800 175.400 153.100 ;
        RECT 179.000 153.100 179.400 153.200 ;
        RECT 179.800 153.100 180.200 153.200 ;
        RECT 179.000 152.800 180.200 153.100 ;
        RECT 59.800 152.100 60.200 152.200 ;
        RECT 65.400 152.100 65.800 152.200 ;
        RECT 59.800 151.800 65.800 152.100 ;
        RECT 109.400 152.100 109.800 152.200 ;
        RECT 111.000 152.100 111.400 152.200 ;
        RECT 119.000 152.100 119.400 152.200 ;
        RECT 109.400 151.800 119.400 152.100 ;
        RECT 123.000 152.100 123.400 152.200 ;
        RECT 143.800 152.100 144.200 152.200 ;
        RECT 146.200 152.100 146.600 152.200 ;
        RECT 123.000 151.800 136.100 152.100 ;
        RECT 143.800 151.800 146.600 152.100 ;
        RECT 167.800 152.100 168.200 152.200 ;
        RECT 183.800 152.100 184.200 152.200 ;
        RECT 167.800 151.800 184.200 152.100 ;
        RECT 135.800 151.200 136.100 151.800 ;
        RECT 11.000 151.100 11.400 151.200 ;
        RECT 61.400 151.100 61.800 151.200 ;
        RECT 11.000 150.800 61.800 151.100 ;
        RECT 67.000 151.100 67.400 151.200 ;
        RECT 69.400 151.100 69.800 151.200 ;
        RECT 67.000 150.800 69.800 151.100 ;
        RECT 75.000 150.800 75.400 151.200 ;
        RECT 107.000 151.100 107.400 151.200 ;
        RECT 119.800 151.100 120.200 151.200 ;
        RECT 123.800 151.100 124.200 151.200 ;
        RECT 107.000 150.800 124.200 151.100 ;
        RECT 128.600 151.100 129.000 151.200 ;
        RECT 133.400 151.100 133.800 151.200 ;
        RECT 128.600 150.800 133.800 151.100 ;
        RECT 135.800 150.800 136.200 151.200 ;
        RECT 177.400 151.100 177.800 151.200 ;
        RECT 184.600 151.100 185.000 151.200 ;
        RECT 177.400 150.800 185.000 151.100 ;
        RECT 194.200 151.100 194.600 151.200 ;
        RECT 196.600 151.100 197.000 151.200 ;
        RECT 194.200 150.800 197.000 151.100 ;
        RECT 75.000 150.200 75.300 150.800 ;
        RECT 15.000 150.100 15.400 150.200 ;
        RECT 39.000 150.100 39.400 150.200 ;
        RECT 15.000 149.800 39.400 150.100 ;
        RECT 55.800 150.100 56.200 150.200 ;
        RECT 71.800 150.100 72.200 150.200 ;
        RECT 55.800 149.800 72.200 150.100 ;
        RECT 75.000 149.800 75.400 150.200 ;
        RECT 111.800 150.100 112.200 150.200 ;
        RECT 124.600 150.100 125.000 150.200 ;
        RECT 125.400 150.100 125.800 150.200 ;
        RECT 111.800 149.800 125.800 150.100 ;
        RECT 135.000 150.100 135.400 150.200 ;
        RECT 140.600 150.100 141.000 150.200 ;
        RECT 135.000 149.800 141.000 150.100 ;
        RECT 159.800 150.100 160.200 150.200 ;
        RECT 163.000 150.100 163.400 150.200 ;
        RECT 178.200 150.100 178.600 150.200 ;
        RECT 159.800 149.800 178.600 150.100 ;
        RECT 182.200 150.100 182.600 150.200 ;
        RECT 183.000 150.100 183.400 150.200 ;
        RECT 182.200 149.800 183.400 150.100 ;
        RECT 183.800 150.100 184.200 150.200 ;
        RECT 191.800 150.100 192.200 150.200 ;
        RECT 183.800 149.800 192.200 150.100 ;
        RECT 10.200 149.100 10.600 149.200 ;
        RECT 14.200 149.100 14.600 149.200 ;
        RECT 10.200 148.800 14.600 149.100 ;
        RECT 27.800 149.100 28.200 149.200 ;
        RECT 62.200 149.100 62.600 149.200 ;
        RECT 27.800 148.800 62.600 149.100 ;
        RECT 63.000 148.800 63.400 149.200 ;
        RECT 75.800 148.800 76.200 149.200 ;
        RECT 86.200 149.100 86.600 149.200 ;
        RECT 95.000 149.100 95.400 149.200 ;
        RECT 86.200 148.800 95.400 149.100 ;
        RECT 125.400 149.100 125.800 149.200 ;
        RECT 143.000 149.100 143.400 149.200 ;
        RECT 125.400 148.800 143.400 149.100 ;
        RECT 152.600 149.100 153.000 149.200 ;
        RECT 154.200 149.100 154.600 149.200 ;
        RECT 152.600 148.800 154.600 149.100 ;
        RECT 169.400 149.100 169.800 149.200 ;
        RECT 170.200 149.100 170.600 149.200 ;
        RECT 169.400 148.800 170.600 149.100 ;
        RECT 171.000 149.100 171.400 149.200 ;
        RECT 173.400 149.100 173.800 149.200 ;
        RECT 171.000 148.800 173.800 149.100 ;
        RECT 174.200 149.100 174.600 149.200 ;
        RECT 181.400 149.100 181.800 149.200 ;
        RECT 191.000 149.100 191.400 149.200 ;
        RECT 174.200 148.800 191.400 149.100 ;
        RECT 63.000 148.200 63.300 148.800 ;
        RECT 9.400 148.100 9.800 148.200 ;
        RECT 16.600 148.100 17.000 148.200 ;
        RECT 25.400 148.100 25.800 148.200 ;
        RECT 9.400 147.800 25.800 148.100 ;
        RECT 26.200 148.100 26.600 148.200 ;
        RECT 35.800 148.100 36.200 148.200 ;
        RECT 26.200 147.800 36.200 148.100 ;
        RECT 49.400 148.100 49.800 148.200 ;
        RECT 54.200 148.100 54.600 148.200 ;
        RECT 55.000 148.100 55.400 148.200 ;
        RECT 49.400 147.800 55.400 148.100 ;
        RECT 63.000 147.800 63.400 148.200 ;
        RECT 66.200 148.100 66.600 148.200 ;
        RECT 75.800 148.100 76.100 148.800 ;
        RECT 66.200 147.800 76.100 148.100 ;
        RECT 83.800 148.100 84.200 148.200 ;
        RECT 84.600 148.100 85.000 148.200 ;
        RECT 83.800 147.800 85.000 148.100 ;
        RECT 119.000 148.100 119.400 148.200 ;
        RECT 120.600 148.100 121.000 148.200 ;
        RECT 119.000 147.800 121.000 148.100 ;
        RECT 121.400 148.100 121.800 148.200 ;
        RECT 131.000 148.100 131.400 148.200 ;
        RECT 121.400 147.800 131.400 148.100 ;
        RECT 146.200 148.100 146.600 148.200 ;
        RECT 151.800 148.100 152.200 148.200 ;
        RECT 161.400 148.100 161.800 148.200 ;
        RECT 167.800 148.100 168.200 148.200 ;
        RECT 146.200 147.800 168.200 148.100 ;
        RECT 168.600 148.100 169.000 148.200 ;
        RECT 174.200 148.100 174.600 148.200 ;
        RECT 168.600 147.800 174.600 148.100 ;
        RECT 177.400 147.800 177.800 148.200 ;
        RECT 182.200 147.800 182.600 148.200 ;
        RECT 183.000 148.100 183.400 148.200 ;
        RECT 184.600 148.100 185.000 148.200 ;
        RECT 183.000 147.800 185.000 148.100 ;
        RECT 195.000 148.100 195.400 148.200 ;
        RECT 202.200 148.100 202.600 148.200 ;
        RECT 195.000 147.800 202.600 148.100 ;
        RECT 3.800 147.100 4.200 147.200 ;
        RECT 11.000 147.100 11.400 147.200 ;
        RECT 12.600 147.100 13.000 147.200 ;
        RECT 17.400 147.100 17.800 147.200 ;
        RECT 3.800 146.800 12.100 147.100 ;
        RECT 12.600 146.800 17.800 147.100 ;
        RECT 19.000 147.100 19.400 147.200 ;
        RECT 24.600 147.100 25.000 147.200 ;
        RECT 19.000 146.800 25.000 147.100 ;
        RECT 35.800 147.100 36.100 147.800 ;
        RECT 44.600 147.100 45.000 147.200 ;
        RECT 35.800 146.800 45.000 147.100 ;
        RECT 46.200 147.100 46.600 147.200 ;
        RECT 55.800 147.100 56.200 147.200 ;
        RECT 46.200 146.800 56.200 147.100 ;
        RECT 57.400 147.100 57.800 147.200 ;
        RECT 58.200 147.100 58.600 147.200 ;
        RECT 57.400 146.800 58.600 147.100 ;
        RECT 63.800 147.100 64.200 147.200 ;
        RECT 86.200 147.100 86.600 147.200 ;
        RECT 63.800 146.800 86.600 147.100 ;
        RECT 89.400 147.100 89.800 147.200 ;
        RECT 95.800 147.100 96.200 147.200 ;
        RECT 89.400 146.800 96.200 147.100 ;
        RECT 104.600 147.100 105.000 147.200 ;
        RECT 111.800 147.100 112.200 147.200 ;
        RECT 104.600 146.800 112.200 147.100 ;
        RECT 118.200 147.100 118.600 147.200 ;
        RECT 123.800 147.100 124.200 147.200 ;
        RECT 118.200 146.800 124.200 147.100 ;
        RECT 137.400 147.100 137.800 147.200 ;
        RECT 174.200 147.100 174.600 147.200 ;
        RECT 137.400 146.800 174.600 147.100 ;
        RECT 177.400 147.100 177.700 147.800 ;
        RECT 182.200 147.100 182.500 147.800 ;
        RECT 187.800 147.100 188.200 147.200 ;
        RECT 194.200 147.100 194.600 147.200 ;
        RECT 197.400 147.100 197.800 147.200 ;
        RECT 177.400 146.800 180.100 147.100 ;
        RECT 182.200 146.800 197.800 147.100 ;
        RECT 11.800 146.100 12.200 146.200 ;
        RECT 14.200 146.100 14.600 146.200 ;
        RECT 18.200 146.100 18.600 146.200 ;
        RECT 24.600 146.100 25.000 146.200 ;
        RECT 11.800 145.800 25.000 146.100 ;
        RECT 51.800 146.100 52.200 146.200 ;
        RECT 54.200 146.100 54.600 146.200 ;
        RECT 51.800 145.800 54.600 146.100 ;
        RECT 99.800 146.100 100.200 146.200 ;
        RECT 103.800 146.100 104.200 146.200 ;
        RECT 99.800 145.800 104.200 146.100 ;
        RECT 106.200 146.100 106.600 146.200 ;
        RECT 122.200 146.100 122.600 146.200 ;
        RECT 129.400 146.100 129.800 146.200 ;
        RECT 131.800 146.100 132.200 146.200 ;
        RECT 136.600 146.100 137.000 146.200 ;
        RECT 143.800 146.100 144.200 146.200 ;
        RECT 155.000 146.100 155.400 146.200 ;
        RECT 157.400 146.100 157.800 146.200 ;
        RECT 179.000 146.100 179.400 146.200 ;
        RECT 106.200 145.800 127.300 146.100 ;
        RECT 129.400 145.800 179.400 146.100 ;
        RECT 179.800 146.100 180.100 146.800 ;
        RECT 185.400 146.100 185.800 146.200 ;
        RECT 179.800 145.800 185.800 146.100 ;
        RECT 187.000 146.100 187.400 146.200 ;
        RECT 187.800 146.100 188.200 146.200 ;
        RECT 187.000 145.800 188.200 146.100 ;
        RECT 127.000 145.200 127.300 145.800 ;
        RECT 12.600 145.100 13.000 145.200 ;
        RECT 13.400 145.100 13.800 145.200 ;
        RECT 21.400 145.100 21.800 145.200 ;
        RECT 12.600 144.800 21.800 145.100 ;
        RECT 51.800 145.100 52.200 145.200 ;
        RECT 54.200 145.100 54.600 145.200 ;
        RECT 51.800 144.800 54.600 145.100 ;
        RECT 59.800 145.100 60.200 145.200 ;
        RECT 102.200 145.100 102.600 145.200 ;
        RECT 105.400 145.100 105.800 145.200 ;
        RECT 59.800 144.800 105.800 145.100 ;
        RECT 115.000 145.100 115.400 145.200 ;
        RECT 117.400 145.100 117.800 145.200 ;
        RECT 115.000 144.800 117.800 145.100 ;
        RECT 120.600 145.100 121.000 145.200 ;
        RECT 125.400 145.100 125.800 145.200 ;
        RECT 120.600 144.800 125.800 145.100 ;
        RECT 127.000 144.800 127.400 145.200 ;
        RECT 127.800 145.100 128.200 145.200 ;
        RECT 129.400 145.100 129.800 145.200 ;
        RECT 127.800 144.800 129.800 145.100 ;
        RECT 147.000 145.100 147.400 145.200 ;
        RECT 159.000 145.100 159.400 145.200 ;
        RECT 147.000 144.800 159.400 145.100 ;
        RECT 171.000 145.100 171.400 145.200 ;
        RECT 171.800 145.100 172.200 145.200 ;
        RECT 171.000 144.800 172.200 145.100 ;
        RECT 180.600 144.800 181.000 145.200 ;
        RECT 182.200 145.100 182.600 145.200 ;
        RECT 183.000 145.100 183.400 145.200 ;
        RECT 190.200 145.100 190.600 145.200 ;
        RECT 182.200 144.800 193.700 145.100 ;
        RECT 10.200 144.100 10.600 144.200 ;
        RECT 13.400 144.100 13.800 144.200 ;
        RECT 10.200 143.800 13.800 144.100 ;
        RECT 19.000 144.100 19.400 144.200 ;
        RECT 20.600 144.100 21.000 144.200 ;
        RECT 19.000 143.800 21.000 144.100 ;
        RECT 59.000 144.100 59.400 144.200 ;
        RECT 110.200 144.100 110.600 144.200 ;
        RECT 59.000 143.800 110.600 144.100 ;
        RECT 117.400 144.100 117.800 144.200 ;
        RECT 120.600 144.100 121.000 144.200 ;
        RECT 117.400 143.800 121.000 144.100 ;
        RECT 123.000 144.100 123.400 144.200 ;
        RECT 126.200 144.100 126.600 144.200 ;
        RECT 128.600 144.100 129.000 144.200 ;
        RECT 123.000 143.800 129.000 144.100 ;
        RECT 135.000 144.100 135.400 144.200 ;
        RECT 142.200 144.100 142.600 144.200 ;
        RECT 135.000 143.800 142.600 144.100 ;
        RECT 148.600 144.100 149.000 144.200 ;
        RECT 163.800 144.100 164.200 144.200 ;
        RECT 180.600 144.100 180.900 144.800 ;
        RECT 193.400 144.200 193.700 144.800 ;
        RECT 201.400 144.800 201.800 145.200 ;
        RECT 201.400 144.200 201.700 144.800 ;
        RECT 148.600 143.800 180.900 144.100 ;
        RECT 185.400 144.100 185.800 144.200 ;
        RECT 187.000 144.100 187.400 144.200 ;
        RECT 185.400 143.800 187.400 144.100 ;
        RECT 193.400 143.800 193.800 144.200 ;
        RECT 194.200 144.100 194.600 144.200 ;
        RECT 196.600 144.100 197.000 144.200 ;
        RECT 194.200 143.800 197.000 144.100 ;
        RECT 201.400 143.800 201.800 144.200 ;
        RECT 22.200 143.100 22.600 143.200 ;
        RECT 55.800 143.100 56.200 143.200 ;
        RECT 58.200 143.100 58.600 143.200 ;
        RECT 87.000 143.100 87.400 143.200 ;
        RECT 89.400 143.100 89.800 143.200 ;
        RECT 100.600 143.100 101.000 143.200 ;
        RECT 107.000 143.100 107.400 143.200 ;
        RECT 22.200 142.800 107.400 143.100 ;
        RECT 118.200 143.100 118.600 143.200 ;
        RECT 123.000 143.100 123.400 143.200 ;
        RECT 124.600 143.100 125.000 143.200 ;
        RECT 127.000 143.100 127.400 143.200 ;
        RECT 118.200 142.800 127.400 143.100 ;
        RECT 127.800 143.100 128.200 143.200 ;
        RECT 145.400 143.100 145.800 143.200 ;
        RECT 175.000 143.100 175.400 143.200 ;
        RECT 127.800 142.800 175.400 143.100 ;
        RECT 191.000 143.100 191.400 143.200 ;
        RECT 195.000 143.100 195.400 143.200 ;
        RECT 191.000 142.800 195.400 143.100 ;
        RECT 199.000 143.100 199.400 143.200 ;
        RECT 199.800 143.100 200.200 143.200 ;
        RECT 199.000 142.800 200.200 143.100 ;
        RECT 19.800 142.100 20.200 142.200 ;
        RECT 30.200 142.100 30.600 142.200 ;
        RECT 19.800 141.800 30.600 142.100 ;
        RECT 67.800 141.800 68.200 142.200 ;
        RECT 115.800 142.100 116.200 142.200 ;
        RECT 138.200 142.100 138.600 142.200 ;
        RECT 145.400 142.100 145.800 142.200 ;
        RECT 115.800 141.800 145.800 142.100 ;
        RECT 149.400 142.100 149.800 142.200 ;
        RECT 161.400 142.100 161.800 142.200 ;
        RECT 149.400 141.800 161.800 142.100 ;
        RECT 167.000 142.100 167.400 142.200 ;
        RECT 171.000 142.100 171.400 142.200 ;
        RECT 191.000 142.100 191.400 142.200 ;
        RECT 167.000 141.800 191.400 142.100 ;
        RECT 192.600 142.100 193.000 142.200 ;
        RECT 195.800 142.100 196.200 142.200 ;
        RECT 192.600 141.800 196.200 142.100 ;
        RECT 67.800 141.200 68.100 141.800 ;
        RECT 67.800 140.800 68.200 141.200 ;
        RECT 92.600 141.100 93.000 141.200 ;
        RECT 118.200 141.100 118.600 141.200 ;
        RECT 92.600 140.800 118.600 141.100 ;
        RECT 123.000 141.100 123.400 141.200 ;
        RECT 128.600 141.100 129.000 141.200 ;
        RECT 123.000 140.800 129.000 141.100 ;
        RECT 131.000 141.100 131.400 141.200 ;
        RECT 147.000 141.100 147.400 141.200 ;
        RECT 131.000 140.800 147.400 141.100 ;
        RECT 155.800 141.100 156.200 141.200 ;
        RECT 171.800 141.100 172.200 141.200 ;
        RECT 155.800 140.800 172.200 141.100 ;
        RECT 172.600 141.100 173.000 141.200 ;
        RECT 173.400 141.100 173.800 141.200 ;
        RECT 172.600 140.800 173.800 141.100 ;
        RECT 176.600 141.100 177.000 141.200 ;
        RECT 199.800 141.100 200.200 141.200 ;
        RECT 176.600 140.800 200.200 141.100 ;
        RECT 78.200 140.100 78.600 140.200 ;
        RECT 80.600 140.100 81.000 140.200 ;
        RECT 103.800 140.100 104.200 140.200 ;
        RECT 107.800 140.100 108.200 140.200 ;
        RECT 115.800 140.100 116.200 140.200 ;
        RECT 141.400 140.100 141.800 140.200 ;
        RECT 78.200 139.800 141.800 140.100 ;
        RECT 172.600 140.100 173.000 140.200 ;
        RECT 173.400 140.100 173.800 140.200 ;
        RECT 172.600 139.800 173.800 140.100 ;
        RECT 183.000 140.100 183.400 140.200 ;
        RECT 192.600 140.100 193.000 140.200 ;
        RECT 183.000 139.800 193.000 140.100 ;
        RECT 20.600 139.100 21.000 139.200 ;
        RECT 21.400 139.100 21.800 139.200 ;
        RECT 20.600 138.800 21.800 139.100 ;
        RECT 107.800 139.100 108.200 139.200 ;
        RECT 109.400 139.100 109.800 139.200 ;
        RECT 127.800 139.100 128.200 139.200 ;
        RECT 107.800 138.800 109.800 139.100 ;
        RECT 110.200 138.800 128.200 139.100 ;
        RECT 128.600 139.100 129.000 139.200 ;
        RECT 148.600 139.100 149.000 139.200 ;
        RECT 128.600 138.800 149.000 139.100 ;
        RECT 155.000 139.100 155.400 139.200 ;
        RECT 155.000 138.800 176.100 139.100 ;
        RECT 70.200 138.100 70.600 138.200 ;
        RECT 103.800 138.100 104.200 138.200 ;
        RECT 70.200 137.800 104.200 138.100 ;
        RECT 105.400 138.100 105.800 138.200 ;
        RECT 110.200 138.100 110.500 138.800 ;
        RECT 175.800 138.200 176.100 138.800 ;
        RECT 105.400 137.800 110.500 138.100 ;
        RECT 111.000 138.100 111.400 138.200 ;
        RECT 113.400 138.100 113.800 138.200 ;
        RECT 127.800 138.100 128.200 138.200 ;
        RECT 140.600 138.100 141.000 138.200 ;
        RECT 111.000 137.800 141.000 138.100 ;
        RECT 161.400 138.100 161.800 138.200 ;
        RECT 170.200 138.100 170.600 138.200 ;
        RECT 172.600 138.100 173.000 138.200 ;
        RECT 161.400 137.800 173.000 138.100 ;
        RECT 175.800 137.800 176.200 138.200 ;
        RECT 199.800 138.100 200.200 138.200 ;
        RECT 176.600 137.800 200.200 138.100 ;
        RECT 202.200 138.100 202.600 138.200 ;
        RECT 203.800 138.100 204.200 138.200 ;
        RECT 202.200 137.800 204.200 138.100 ;
        RECT 46.200 137.100 46.600 137.200 ;
        RECT 52.600 137.100 53.000 137.200 ;
        RECT 46.200 136.800 53.000 137.100 ;
        RECT 91.800 136.800 92.200 137.200 ;
        RECT 101.400 137.100 101.800 137.200 ;
        RECT 119.000 137.100 119.400 137.200 ;
        RECT 101.400 136.800 119.400 137.100 ;
        RECT 125.400 136.800 125.800 137.200 ;
        RECT 126.200 137.100 126.600 137.200 ;
        RECT 127.000 137.100 127.400 137.200 ;
        RECT 126.200 136.800 127.400 137.100 ;
        RECT 144.600 137.100 145.000 137.200 ;
        RECT 164.600 137.100 165.000 137.200 ;
        RECT 144.600 136.800 165.000 137.100 ;
        RECT 175.000 137.100 175.400 137.200 ;
        RECT 176.600 137.100 176.900 137.800 ;
        RECT 175.000 136.800 176.900 137.100 ;
        RECT 178.200 137.100 178.600 137.200 ;
        RECT 184.600 137.100 185.000 137.200 ;
        RECT 178.200 136.800 185.000 137.100 ;
        RECT 91.800 136.200 92.100 136.800 ;
        RECT 125.400 136.200 125.700 136.800 ;
        RECT 13.400 136.100 13.800 136.200 ;
        RECT 38.200 136.100 38.600 136.200 ;
        RECT 13.400 135.800 38.600 136.100 ;
        RECT 65.400 135.800 65.800 136.200 ;
        RECT 66.200 135.800 66.600 136.200 ;
        RECT 68.600 136.100 69.000 136.200 ;
        RECT 73.400 136.100 73.800 136.200 ;
        RECT 68.600 135.800 73.800 136.100 ;
        RECT 88.600 135.800 89.000 136.200 ;
        RECT 91.800 135.800 92.200 136.200 ;
        RECT 95.800 136.100 96.200 136.200 ;
        RECT 102.200 136.100 102.600 136.200 ;
        RECT 120.600 136.100 121.000 136.200 ;
        RECT 95.800 135.800 121.000 136.100 ;
        RECT 125.400 135.800 125.800 136.200 ;
        RECT 131.800 136.100 132.200 136.200 ;
        RECT 134.200 136.100 134.600 136.200 ;
        RECT 149.400 136.100 149.800 136.200 ;
        RECT 161.400 136.100 161.800 136.200 ;
        RECT 131.800 135.800 134.600 136.100 ;
        RECT 148.600 135.800 161.800 136.100 ;
        RECT 166.200 135.800 166.600 136.200 ;
        RECT 179.000 136.100 179.400 136.200 ;
        RECT 180.600 136.100 181.000 136.200 ;
        RECT 179.000 135.800 181.000 136.100 ;
        RECT 187.800 136.100 188.200 136.200 ;
        RECT 189.400 136.100 189.800 136.200 ;
        RECT 193.400 136.100 193.800 136.200 ;
        RECT 187.800 135.800 193.800 136.100 ;
        RECT 195.800 136.100 196.200 136.200 ;
        RECT 197.400 136.100 197.800 136.200 ;
        RECT 195.800 135.800 197.800 136.100 ;
        RECT 198.200 136.100 198.600 136.200 ;
        RECT 199.000 136.100 199.400 136.200 ;
        RECT 198.200 135.800 199.400 136.100 ;
        RECT 18.200 135.100 18.600 135.200 ;
        RECT 19.000 135.100 19.400 135.200 ;
        RECT 18.200 134.800 19.400 135.100 ;
        RECT 42.200 135.100 42.600 135.200 ;
        RECT 47.000 135.100 47.400 135.200 ;
        RECT 49.400 135.100 49.800 135.200 ;
        RECT 42.200 134.800 49.800 135.100 ;
        RECT 56.600 135.100 57.000 135.200 ;
        RECT 65.400 135.100 65.700 135.800 ;
        RECT 56.600 134.800 65.700 135.100 ;
        RECT 66.200 135.200 66.500 135.800 ;
        RECT 66.200 134.800 66.600 135.200 ;
        RECT 70.200 135.100 70.600 135.200 ;
        RECT 74.200 135.100 74.600 135.200 ;
        RECT 70.200 134.800 74.600 135.100 ;
        RECT 77.400 135.100 77.800 135.200 ;
        RECT 79.000 135.100 79.400 135.200 ;
        RECT 77.400 134.800 79.400 135.100 ;
        RECT 88.600 135.100 88.900 135.800 ;
        RECT 94.200 135.100 94.600 135.200 ;
        RECT 88.600 134.800 94.600 135.100 ;
        RECT 109.400 135.100 109.800 135.200 ;
        RECT 114.200 135.100 114.600 135.200 ;
        RECT 123.000 135.100 123.400 135.200 ;
        RECT 109.400 134.800 114.600 135.100 ;
        RECT 121.400 134.800 123.400 135.100 ;
        RECT 131.000 135.100 131.400 135.200 ;
        RECT 135.800 135.100 136.200 135.200 ;
        RECT 131.000 134.800 136.200 135.100 ;
        RECT 137.400 135.100 137.800 135.200 ;
        RECT 138.200 135.100 138.600 135.200 ;
        RECT 137.400 134.800 138.600 135.100 ;
        RECT 142.200 135.100 142.600 135.200 ;
        RECT 146.200 135.100 146.600 135.200 ;
        RECT 142.200 134.800 146.600 135.100 ;
        RECT 152.600 134.800 153.000 135.200 ;
        RECT 164.600 135.100 165.000 135.200 ;
        RECT 166.200 135.100 166.500 135.800 ;
        RECT 164.600 134.800 166.500 135.100 ;
        RECT 173.400 135.100 173.800 135.200 ;
        RECT 178.200 135.100 178.600 135.200 ;
        RECT 179.800 135.100 180.200 135.200 ;
        RECT 183.800 135.100 184.200 135.200 ;
        RECT 173.400 134.800 179.300 135.100 ;
        RECT 179.800 134.800 197.700 135.100 ;
        RECT 121.400 134.700 121.800 134.800 ;
        RECT 9.400 133.800 9.800 134.200 ;
        RECT 15.800 134.100 16.200 134.200 ;
        RECT 25.400 134.100 25.800 134.200 ;
        RECT 15.800 133.800 25.800 134.100 ;
        RECT 39.000 134.100 39.400 134.200 ;
        RECT 41.400 134.100 41.800 134.200 ;
        RECT 39.000 133.800 41.800 134.100 ;
        RECT 47.800 133.800 48.200 134.200 ;
        RECT 52.600 134.100 53.000 134.200 ;
        RECT 63.800 134.100 64.200 134.200 ;
        RECT 66.200 134.100 66.600 134.200 ;
        RECT 69.400 134.100 69.800 134.200 ;
        RECT 71.000 134.100 71.400 134.200 ;
        RECT 93.400 134.100 93.800 134.200 ;
        RECT 97.400 134.100 97.800 134.200 ;
        RECT 128.600 134.100 129.000 134.200 ;
        RECT 52.600 133.800 129.000 134.100 ;
        RECT 136.600 134.100 137.000 134.200 ;
        RECT 138.200 134.100 138.600 134.200 ;
        RECT 136.600 133.800 138.600 134.100 ;
        RECT 151.800 134.100 152.200 134.200 ;
        RECT 152.600 134.100 152.900 134.800 ;
        RECT 197.400 134.200 197.700 134.800 ;
        RECT 151.800 133.800 152.900 134.100 ;
        RECT 167.800 134.100 168.200 134.200 ;
        RECT 178.200 134.100 178.600 134.200 ;
        RECT 179.000 134.100 179.400 134.200 ;
        RECT 167.800 133.800 179.400 134.100 ;
        RECT 179.800 134.100 180.200 134.200 ;
        RECT 186.200 134.100 186.600 134.200 ;
        RECT 179.800 133.800 186.600 134.100 ;
        RECT 192.600 134.100 193.000 134.200 ;
        RECT 194.200 134.100 194.600 134.200 ;
        RECT 196.600 134.100 197.000 134.200 ;
        RECT 192.600 133.800 197.000 134.100 ;
        RECT 197.400 134.100 197.800 134.200 ;
        RECT 198.200 134.100 198.600 134.200 ;
        RECT 197.400 133.800 198.600 134.100 ;
        RECT 3.000 133.100 3.400 133.200 ;
        RECT 9.400 133.100 9.700 133.800 ;
        RECT 23.000 133.100 23.400 133.200 ;
        RECT 40.600 133.100 41.000 133.200 ;
        RECT 42.200 133.100 42.600 133.200 ;
        RECT 3.000 132.800 29.700 133.100 ;
        RECT 40.600 132.800 42.600 133.100 ;
        RECT 45.400 133.100 45.800 133.200 ;
        RECT 47.800 133.100 48.100 133.800 ;
        RECT 45.400 132.800 48.100 133.100 ;
        RECT 55.800 133.100 56.200 133.200 ;
        RECT 80.600 133.100 81.000 133.200 ;
        RECT 125.400 133.100 125.800 133.200 ;
        RECT 131.800 133.100 132.200 133.200 ;
        RECT 55.800 132.800 98.500 133.100 ;
        RECT 125.400 132.800 132.200 133.100 ;
        RECT 134.200 133.100 134.600 133.200 ;
        RECT 165.400 133.100 165.800 133.200 ;
        RECT 134.200 132.800 165.800 133.100 ;
        RECT 181.400 133.100 181.800 133.200 ;
        RECT 183.800 133.100 184.200 133.200 ;
        RECT 200.600 133.100 201.000 133.200 ;
        RECT 181.400 132.800 201.000 133.100 ;
        RECT 29.400 132.200 29.700 132.800 ;
        RECT 98.200 132.200 98.500 132.800 ;
        RECT 29.400 131.800 29.800 132.200 ;
        RECT 39.800 132.100 40.200 132.200 ;
        RECT 44.600 132.100 45.000 132.200 ;
        RECT 39.800 131.800 45.000 132.100 ;
        RECT 52.600 132.100 53.000 132.200 ;
        RECT 59.800 132.100 60.200 132.200 ;
        RECT 52.600 131.800 60.200 132.100 ;
        RECT 67.000 132.100 67.400 132.200 ;
        RECT 67.800 132.100 68.200 132.200 ;
        RECT 75.800 132.100 76.200 132.200 ;
        RECT 80.600 132.100 81.000 132.200 ;
        RECT 67.000 131.800 81.000 132.100 ;
        RECT 81.400 132.100 81.800 132.200 ;
        RECT 82.200 132.100 82.600 132.200 ;
        RECT 81.400 131.800 82.600 132.100 ;
        RECT 98.200 131.800 98.600 132.200 ;
        RECT 99.800 132.100 100.200 132.200 ;
        RECT 107.800 132.100 108.200 132.200 ;
        RECT 99.800 131.800 108.200 132.100 ;
        RECT 110.200 132.100 110.600 132.200 ;
        RECT 135.800 132.100 136.200 132.200 ;
        RECT 110.200 131.800 136.200 132.100 ;
        RECT 156.600 132.100 157.000 132.200 ;
        RECT 167.000 132.100 167.400 132.200 ;
        RECT 156.600 131.800 167.400 132.100 ;
        RECT 176.600 132.100 177.000 132.200 ;
        RECT 179.800 132.100 180.200 132.200 ;
        RECT 176.600 131.800 180.200 132.100 ;
        RECT 186.200 132.100 186.600 132.200 ;
        RECT 195.800 132.100 196.200 132.200 ;
        RECT 186.200 131.800 196.200 132.100 ;
        RECT 11.000 131.100 11.400 131.200 ;
        RECT 41.400 131.100 41.800 131.200 ;
        RECT 11.000 130.800 41.800 131.100 ;
        RECT 43.000 131.100 43.400 131.200 ;
        RECT 43.800 131.100 44.200 131.200 ;
        RECT 43.000 130.800 44.200 131.100 ;
        RECT 44.600 131.100 45.000 131.200 ;
        RECT 55.800 131.100 56.200 131.200 ;
        RECT 44.600 130.800 56.200 131.100 ;
        RECT 75.800 131.100 76.200 131.200 ;
        RECT 76.600 131.100 77.000 131.200 ;
        RECT 75.800 130.800 77.000 131.100 ;
        RECT 78.200 131.100 78.600 131.200 ;
        RECT 87.000 131.100 87.400 131.200 ;
        RECT 92.600 131.100 93.000 131.200 ;
        RECT 78.200 130.800 93.000 131.100 ;
        RECT 104.600 131.100 105.000 131.200 ;
        RECT 115.000 131.100 115.400 131.200 ;
        RECT 104.600 130.800 115.400 131.100 ;
        RECT 115.800 131.100 116.200 131.200 ;
        RECT 117.400 131.100 117.800 131.200 ;
        RECT 135.000 131.100 135.400 131.200 ;
        RECT 115.800 130.800 135.400 131.100 ;
        RECT 146.200 131.100 146.600 131.200 ;
        RECT 171.000 131.100 171.400 131.200 ;
        RECT 146.200 130.800 171.400 131.100 ;
        RECT 15.000 130.100 15.400 130.200 ;
        RECT 44.600 130.100 45.000 130.200 ;
        RECT 15.000 129.800 45.000 130.100 ;
        RECT 49.400 129.800 49.800 130.200 ;
        RECT 82.200 130.100 82.600 130.200 ;
        RECT 87.000 130.100 87.400 130.200 ;
        RECT 91.800 130.100 92.200 130.200 ;
        RECT 82.200 129.800 92.200 130.100 ;
        RECT 115.000 130.100 115.400 130.200 ;
        RECT 118.200 130.100 118.600 130.200 ;
        RECT 115.000 129.800 118.600 130.100 ;
        RECT 139.800 130.100 140.200 130.200 ;
        RECT 160.600 130.100 161.000 130.200 ;
        RECT 168.600 130.100 169.000 130.200 ;
        RECT 187.000 130.100 187.400 130.200 ;
        RECT 139.800 129.800 187.400 130.100 ;
        RECT 189.400 130.100 189.800 130.200 ;
        RECT 195.000 130.100 195.400 130.200 ;
        RECT 196.600 130.100 197.000 130.200 ;
        RECT 189.400 129.800 197.000 130.100 ;
        RECT 198.200 130.100 198.600 130.200 ;
        RECT 199.000 130.100 199.400 130.200 ;
        RECT 198.200 129.800 199.400 130.100 ;
        RECT 199.800 130.100 200.200 130.200 ;
        RECT 203.000 130.100 203.400 130.200 ;
        RECT 199.800 129.800 203.400 130.100 ;
        RECT 11.000 128.800 11.400 129.200 ;
        RECT 27.000 129.100 27.400 129.200 ;
        RECT 29.400 129.100 29.800 129.200 ;
        RECT 39.000 129.100 39.400 129.200 ;
        RECT 43.000 129.100 43.400 129.200 ;
        RECT 27.000 128.800 43.400 129.100 ;
        RECT 43.800 129.100 44.200 129.200 ;
        RECT 45.400 129.100 45.800 129.200 ;
        RECT 48.600 129.100 49.000 129.200 ;
        RECT 49.400 129.100 49.700 129.800 ;
        RECT 43.800 128.800 46.500 129.100 ;
        RECT 48.600 128.800 49.700 129.100 ;
        RECT 50.200 129.100 50.600 129.200 ;
        RECT 57.400 129.100 57.800 129.200 ;
        RECT 50.200 128.800 57.800 129.100 ;
        RECT 70.200 129.100 70.600 129.200 ;
        RECT 89.400 129.100 89.800 129.200 ;
        RECT 70.200 128.800 89.800 129.100 ;
        RECT 90.200 129.100 90.600 129.200 ;
        RECT 99.000 129.100 99.400 129.200 ;
        RECT 90.200 128.800 99.400 129.100 ;
        RECT 109.400 128.800 109.800 129.200 ;
        RECT 115.800 128.800 116.200 129.200 ;
        RECT 137.400 129.100 137.800 129.200 ;
        RECT 142.200 129.100 142.600 129.200 ;
        RECT 137.400 128.800 142.600 129.100 ;
        RECT 145.400 129.100 145.800 129.200 ;
        RECT 154.200 129.100 154.600 129.200 ;
        RECT 145.400 128.800 154.600 129.100 ;
        RECT 155.800 129.100 156.200 129.200 ;
        RECT 175.800 129.100 176.200 129.200 ;
        RECT 176.600 129.100 177.000 129.200 ;
        RECT 155.800 128.800 169.700 129.100 ;
        RECT 175.800 128.800 177.000 129.100 ;
        RECT 183.800 129.100 184.200 129.200 ;
        RECT 187.800 129.100 188.200 129.200 ;
        RECT 183.800 128.800 188.200 129.100 ;
        RECT 11.000 128.100 11.300 128.800 ;
        RECT 109.400 128.200 109.700 128.800 ;
        RECT 115.800 128.200 116.100 128.800 ;
        RECT 169.400 128.200 169.700 128.800 ;
        RECT 15.000 128.100 15.400 128.200 ;
        RECT 11.000 127.800 15.400 128.100 ;
        RECT 19.800 128.100 20.200 128.200 ;
        RECT 28.600 128.100 29.000 128.200 ;
        RECT 19.800 127.800 29.000 128.100 ;
        RECT 31.000 128.100 31.400 128.200 ;
        RECT 40.600 128.100 41.000 128.200 ;
        RECT 31.000 127.800 41.000 128.100 ;
        RECT 43.800 128.100 44.200 128.200 ;
        RECT 47.000 128.100 47.400 128.200 ;
        RECT 43.800 127.800 47.400 128.100 ;
        RECT 50.200 128.100 50.600 128.200 ;
        RECT 59.800 128.100 60.200 128.200 ;
        RECT 50.200 127.800 60.200 128.100 ;
        RECT 60.600 128.100 61.000 128.200 ;
        RECT 67.800 128.100 68.200 128.200 ;
        RECT 60.600 127.800 68.200 128.100 ;
        RECT 83.000 128.100 83.400 128.200 ;
        RECT 83.800 128.100 84.200 128.200 ;
        RECT 83.000 127.800 84.200 128.100 ;
        RECT 84.600 128.100 85.000 128.200 ;
        RECT 85.400 128.100 85.800 128.200 ;
        RECT 84.600 127.800 85.800 128.100 ;
        RECT 87.000 128.100 87.400 128.200 ;
        RECT 88.600 128.100 89.000 128.200 ;
        RECT 87.000 127.800 89.000 128.100 ;
        RECT 108.600 127.800 109.000 128.200 ;
        RECT 109.400 127.800 109.800 128.200 ;
        RECT 115.800 127.800 116.200 128.200 ;
        RECT 131.000 128.100 131.400 128.200 ;
        RECT 139.000 128.100 139.400 128.200 ;
        RECT 131.000 127.800 139.400 128.100 ;
        RECT 162.200 128.100 162.600 128.200 ;
        RECT 162.200 127.800 164.900 128.100 ;
        RECT 169.400 127.800 169.800 128.200 ;
        RECT 171.000 128.100 171.400 128.200 ;
        RECT 174.200 128.100 174.600 128.200 ;
        RECT 171.000 127.800 174.600 128.100 ;
        RECT 177.400 128.100 177.800 128.200 ;
        RECT 179.800 128.100 180.200 128.200 ;
        RECT 183.800 128.100 184.100 128.800 ;
        RECT 193.400 128.100 193.800 128.200 ;
        RECT 177.400 127.800 184.100 128.100 ;
        RECT 187.000 127.800 193.800 128.100 ;
        RECT 202.200 128.100 202.600 128.200 ;
        RECT 203.000 128.100 203.400 128.200 ;
        RECT 202.200 127.800 203.400 128.100 ;
        RECT 5.400 127.100 5.800 127.200 ;
        RECT 11.800 127.100 12.200 127.200 ;
        RECT 5.400 126.800 12.200 127.100 ;
        RECT 25.400 127.100 25.800 127.200 ;
        RECT 31.000 127.100 31.400 127.200 ;
        RECT 47.000 127.100 47.400 127.200 ;
        RECT 47.800 127.100 48.200 127.200 ;
        RECT 25.400 126.800 42.500 127.100 ;
        RECT 47.000 126.800 48.200 127.100 ;
        RECT 48.600 127.100 49.000 127.200 ;
        RECT 58.200 127.100 58.600 127.200 ;
        RECT 59.000 127.100 59.400 127.200 ;
        RECT 48.600 126.800 57.700 127.100 ;
        RECT 58.200 126.800 59.400 127.100 ;
        RECT 66.200 127.100 66.600 127.200 ;
        RECT 67.000 127.100 67.400 127.200 ;
        RECT 66.200 126.800 67.400 127.100 ;
        RECT 70.200 127.100 70.600 127.200 ;
        RECT 86.200 127.100 86.600 127.200 ;
        RECT 103.800 127.100 104.200 127.200 ;
        RECT 104.600 127.100 105.000 127.200 ;
        RECT 70.200 126.800 105.000 127.100 ;
        RECT 106.200 127.100 106.600 127.200 ;
        RECT 107.800 127.100 108.200 127.200 ;
        RECT 106.200 126.800 108.200 127.100 ;
        RECT 108.600 127.100 108.900 127.800 ;
        RECT 164.600 127.200 164.900 127.800 ;
        RECT 110.200 127.100 110.600 127.200 ;
        RECT 108.600 126.800 110.600 127.100 ;
        RECT 138.200 127.100 138.600 127.200 ;
        RECT 139.000 127.100 139.400 127.200 ;
        RECT 138.200 126.800 139.400 127.100 ;
        RECT 151.000 127.100 151.400 127.200 ;
        RECT 157.400 127.100 157.800 127.200 ;
        RECT 151.000 126.800 157.800 127.100 ;
        RECT 159.000 127.100 159.400 127.200 ;
        RECT 162.200 127.100 162.600 127.200 ;
        RECT 159.000 126.800 162.600 127.100 ;
        RECT 164.600 126.800 165.000 127.200 ;
        RECT 168.600 127.100 169.000 127.200 ;
        RECT 169.400 127.100 169.800 127.200 ;
        RECT 168.600 126.800 169.800 127.100 ;
        RECT 172.600 127.100 173.000 127.200 ;
        RECT 187.000 127.100 187.300 127.800 ;
        RECT 172.600 126.800 187.300 127.100 ;
        RECT 187.800 127.100 188.200 127.200 ;
        RECT 195.800 127.100 196.200 127.200 ;
        RECT 187.800 126.800 196.200 127.100 ;
        RECT 201.400 127.100 201.800 127.200 ;
        RECT 203.800 127.100 204.200 127.200 ;
        RECT 201.400 126.800 204.200 127.100 ;
        RECT 12.600 126.100 13.000 126.200 ;
        RECT 13.400 126.100 13.800 126.200 ;
        RECT 21.400 126.100 21.800 126.200 ;
        RECT 12.600 125.800 13.800 126.100 ;
        RECT 15.800 125.800 21.800 126.100 ;
        RECT 24.600 126.100 25.000 126.200 ;
        RECT 26.200 126.100 26.600 126.200 ;
        RECT 34.200 126.100 34.600 126.200 ;
        RECT 35.000 126.100 35.400 126.200 ;
        RECT 24.600 125.800 35.400 126.100 ;
        RECT 36.600 126.100 37.000 126.200 ;
        RECT 40.600 126.100 41.000 126.200 ;
        RECT 36.600 125.800 41.000 126.100 ;
        RECT 42.200 126.100 42.500 126.800 ;
        RECT 51.000 126.100 51.400 126.200 ;
        RECT 42.200 125.800 51.400 126.100 ;
        RECT 57.400 126.100 57.700 126.800 ;
        RECT 66.200 126.100 66.600 126.200 ;
        RECT 76.600 126.100 77.000 126.200 ;
        RECT 57.400 125.800 66.600 126.100 ;
        RECT 71.000 125.800 77.000 126.100 ;
        RECT 80.600 126.100 81.000 126.200 ;
        RECT 86.200 126.100 86.600 126.200 ;
        RECT 80.600 125.800 86.600 126.100 ;
        RECT 94.200 126.100 94.600 126.200 ;
        RECT 99.800 126.100 100.200 126.200 ;
        RECT 94.200 125.800 100.200 126.100 ;
        RECT 100.600 126.100 101.000 126.200 ;
        RECT 105.400 126.100 105.800 126.200 ;
        RECT 111.000 126.100 111.400 126.200 ;
        RECT 100.600 125.800 111.400 126.100 ;
        RECT 112.600 126.100 113.000 126.200 ;
        RECT 123.000 126.100 123.400 126.200 ;
        RECT 112.600 125.800 123.400 126.100 ;
        RECT 139.000 126.100 139.400 126.200 ;
        RECT 139.800 126.100 140.200 126.200 ;
        RECT 140.600 126.100 141.000 126.200 ;
        RECT 139.000 125.800 141.000 126.100 ;
        RECT 158.200 126.100 158.600 126.200 ;
        RECT 159.800 126.100 160.200 126.200 ;
        RECT 158.200 125.800 160.200 126.100 ;
        RECT 161.400 126.100 161.800 126.200 ;
        RECT 162.200 126.100 162.600 126.200 ;
        RECT 161.400 125.800 162.600 126.100 ;
        RECT 163.800 126.100 164.200 126.200 ;
        RECT 167.800 126.100 168.200 126.200 ;
        RECT 173.400 126.100 173.800 126.200 ;
        RECT 163.800 125.800 173.800 126.100 ;
        RECT 174.200 126.100 174.600 126.200 ;
        RECT 191.800 126.100 192.200 126.200 ;
        RECT 194.200 126.100 194.600 126.200 ;
        RECT 199.800 126.100 200.200 126.200 ;
        RECT 174.200 125.800 192.200 126.100 ;
        RECT 193.400 125.800 200.200 126.100 ;
        RECT 15.800 125.200 16.100 125.800 ;
        RECT 71.000 125.200 71.300 125.800 ;
        RECT 15.800 124.800 16.200 125.200 ;
        RECT 19.800 125.100 20.200 125.200 ;
        RECT 27.800 125.100 28.200 125.200 ;
        RECT 19.800 124.800 28.200 125.100 ;
        RECT 37.400 125.100 37.800 125.200 ;
        RECT 54.200 125.100 54.600 125.200 ;
        RECT 67.800 125.100 68.200 125.200 ;
        RECT 37.400 124.800 68.200 125.100 ;
        RECT 71.000 124.800 71.400 125.200 ;
        RECT 75.800 125.100 76.200 125.200 ;
        RECT 83.000 125.100 83.400 125.200 ;
        RECT 75.800 124.800 83.400 125.100 ;
        RECT 107.800 125.100 108.200 125.200 ;
        RECT 131.000 125.100 131.400 125.200 ;
        RECT 107.800 124.800 131.400 125.100 ;
        RECT 135.000 125.100 135.400 125.200 ;
        RECT 142.200 125.100 142.600 125.200 ;
        RECT 147.800 125.100 148.200 125.200 ;
        RECT 135.000 124.800 148.200 125.100 ;
        RECT 165.400 125.100 165.800 125.200 ;
        RECT 171.800 125.100 172.200 125.200 ;
        RECT 165.400 124.800 172.200 125.100 ;
        RECT 174.200 125.100 174.600 125.200 ;
        RECT 182.200 125.100 182.600 125.200 ;
        RECT 183.800 125.100 184.200 125.200 ;
        RECT 174.200 124.800 184.200 125.100 ;
        RECT 37.400 124.200 37.700 124.800 ;
        RECT 171.800 124.200 172.100 124.800 ;
        RECT 37.400 123.800 37.800 124.200 ;
        RECT 43.800 124.100 44.200 124.200 ;
        RECT 46.200 124.100 46.600 124.200 ;
        RECT 43.800 123.800 46.600 124.100 ;
        RECT 53.400 124.100 53.800 124.200 ;
        RECT 55.800 124.100 56.200 124.200 ;
        RECT 65.400 124.100 65.800 124.200 ;
        RECT 74.200 124.100 74.600 124.200 ;
        RECT 84.600 124.100 85.000 124.200 ;
        RECT 53.400 123.800 85.000 124.100 ;
        RECT 86.200 124.100 86.600 124.200 ;
        RECT 113.400 124.100 113.800 124.200 ;
        RECT 86.200 123.800 113.800 124.100 ;
        RECT 116.600 124.100 117.000 124.200 ;
        RECT 122.200 124.100 122.600 124.200 ;
        RECT 116.600 123.800 122.600 124.100 ;
        RECT 165.400 124.100 165.800 124.200 ;
        RECT 171.000 124.100 171.400 124.200 ;
        RECT 165.400 123.800 171.400 124.100 ;
        RECT 171.800 123.800 172.200 124.200 ;
        RECT 172.600 124.100 173.000 124.200 ;
        RECT 174.200 124.100 174.600 124.200 ;
        RECT 172.600 123.800 174.600 124.100 ;
        RECT 198.200 124.100 198.600 124.200 ;
        RECT 204.600 124.100 205.000 124.200 ;
        RECT 198.200 123.800 205.000 124.100 ;
        RECT 44.600 123.100 45.000 123.200 ;
        RECT 47.800 123.100 48.200 123.200 ;
        RECT 44.600 122.800 48.200 123.100 ;
        RECT 49.400 123.100 49.800 123.200 ;
        RECT 53.400 123.100 53.800 123.200 ;
        RECT 63.000 123.100 63.400 123.200 ;
        RECT 49.400 122.800 53.800 123.100 ;
        RECT 55.000 122.800 63.400 123.100 ;
        RECT 67.800 123.100 68.200 123.200 ;
        RECT 78.200 123.100 78.600 123.200 ;
        RECT 67.800 122.800 78.600 123.100 ;
        RECT 79.000 123.100 79.400 123.200 ;
        RECT 106.200 123.100 106.600 123.200 ;
        RECT 79.000 122.800 106.600 123.100 ;
        RECT 110.200 123.100 110.600 123.200 ;
        RECT 117.400 123.100 117.800 123.200 ;
        RECT 110.200 122.800 117.800 123.100 ;
        RECT 163.000 122.800 163.400 123.200 ;
        RECT 55.000 122.200 55.300 122.800 ;
        RECT 163.000 122.200 163.300 122.800 ;
        RECT 43.800 122.100 44.200 122.200 ;
        RECT 47.000 122.100 47.400 122.200 ;
        RECT 43.800 121.800 47.400 122.100 ;
        RECT 55.000 121.800 55.400 122.200 ;
        RECT 75.000 122.100 75.400 122.200 ;
        RECT 76.600 122.100 77.000 122.200 ;
        RECT 75.000 121.800 77.000 122.100 ;
        RECT 111.800 122.100 112.200 122.200 ;
        RECT 123.000 122.100 123.400 122.200 ;
        RECT 111.800 121.800 123.400 122.100 ;
        RECT 163.000 121.800 163.400 122.200 ;
        RECT 188.600 121.800 189.000 122.200 ;
        RECT 191.000 121.800 191.400 122.200 ;
        RECT 188.600 121.200 188.900 121.800 ;
        RECT 191.000 121.200 191.300 121.800 ;
        RECT 68.600 121.100 69.000 121.200 ;
        RECT 81.400 121.100 81.800 121.200 ;
        RECT 68.600 120.800 81.800 121.100 ;
        RECT 159.800 120.800 160.200 121.200 ;
        RECT 163.000 121.100 163.400 121.200 ;
        RECT 173.400 121.100 173.800 121.200 ;
        RECT 163.000 120.800 173.800 121.100 ;
        RECT 188.600 120.800 189.000 121.200 ;
        RECT 191.000 120.800 191.400 121.200 ;
        RECT 159.800 120.200 160.100 120.800 ;
        RECT 123.800 120.100 124.200 120.200 ;
        RECT 144.600 120.100 145.000 120.200 ;
        RECT 123.800 119.800 145.000 120.100 ;
        RECT 159.800 119.800 160.200 120.200 ;
        RECT 61.400 119.100 61.800 119.200 ;
        RECT 63.800 119.100 64.200 119.200 ;
        RECT 61.400 118.800 64.200 119.100 ;
        RECT 83.800 119.100 84.200 119.200 ;
        RECT 107.800 119.100 108.200 119.200 ;
        RECT 83.800 118.800 108.200 119.100 ;
        RECT 108.600 119.100 109.000 119.200 ;
        RECT 170.200 119.100 170.600 119.200 ;
        RECT 108.600 118.800 170.600 119.100 ;
        RECT 183.800 118.800 184.200 119.200 ;
        RECT 39.800 118.100 40.200 118.200 ;
        RECT 46.200 118.100 46.600 118.200 ;
        RECT 39.800 117.800 46.600 118.100 ;
        RECT 58.200 118.100 58.600 118.200 ;
        RECT 63.800 118.100 64.200 118.200 ;
        RECT 64.600 118.100 65.000 118.200 ;
        RECT 58.200 117.800 65.000 118.100 ;
        RECT 85.400 118.100 85.800 118.200 ;
        RECT 86.200 118.100 86.600 118.200 ;
        RECT 85.400 117.800 86.600 118.100 ;
        RECT 87.000 118.100 87.400 118.200 ;
        RECT 149.400 118.100 149.800 118.200 ;
        RECT 167.000 118.100 167.400 118.200 ;
        RECT 183.800 118.100 184.100 118.800 ;
        RECT 87.000 117.800 129.700 118.100 ;
        RECT 149.400 117.800 162.500 118.100 ;
        RECT 167.000 117.800 184.100 118.100 ;
        RECT 129.400 117.200 129.700 117.800 ;
        RECT 43.000 117.100 43.400 117.200 ;
        RECT 58.200 117.100 58.600 117.200 ;
        RECT 91.800 117.100 92.200 117.200 ;
        RECT 43.000 116.800 92.200 117.100 ;
        RECT 119.000 116.800 119.400 117.200 ;
        RECT 129.400 116.800 129.800 117.200 ;
        RECT 132.600 117.100 133.000 117.200 ;
        RECT 151.800 117.100 152.200 117.200 ;
        RECT 132.600 116.800 152.200 117.100 ;
        RECT 162.200 117.100 162.500 117.800 ;
        RECT 169.400 117.100 169.800 117.200 ;
        RECT 162.200 116.800 169.800 117.100 ;
        RECT 22.200 116.100 22.600 116.200 ;
        RECT 42.200 116.100 42.600 116.200 ;
        RECT 22.200 115.800 42.600 116.100 ;
        RECT 53.400 116.100 53.800 116.200 ;
        RECT 65.400 116.100 65.800 116.200 ;
        RECT 86.200 116.100 86.600 116.200 ;
        RECT 53.400 115.800 86.600 116.100 ;
        RECT 87.800 116.100 88.200 116.200 ;
        RECT 91.800 116.100 92.100 116.800 ;
        RECT 119.000 116.200 119.300 116.800 ;
        RECT 92.600 116.100 93.000 116.200 ;
        RECT 87.800 115.800 93.000 116.100 ;
        RECT 96.600 116.100 97.000 116.200 ;
        RECT 106.200 116.100 106.600 116.200 ;
        RECT 96.600 115.800 106.600 116.100 ;
        RECT 109.400 115.800 109.800 116.200 ;
        RECT 119.000 116.100 119.400 116.200 ;
        RECT 120.600 116.100 121.000 116.200 ;
        RECT 119.000 115.800 121.000 116.100 ;
        RECT 138.200 115.800 138.600 116.200 ;
        RECT 143.800 116.100 144.200 116.200 ;
        RECT 145.400 116.100 145.800 116.200 ;
        RECT 143.800 115.800 145.800 116.100 ;
        RECT 151.800 116.100 152.100 116.800 ;
        RECT 157.400 116.100 157.800 116.200 ;
        RECT 159.800 116.100 160.200 116.200 ;
        RECT 163.000 116.100 163.400 116.200 ;
        RECT 151.800 115.800 163.400 116.100 ;
        RECT 164.600 116.100 165.000 116.200 ;
        RECT 166.200 116.100 166.600 116.200 ;
        RECT 164.600 115.800 166.600 116.100 ;
        RECT 175.800 116.100 176.200 116.200 ;
        RECT 202.200 116.100 202.600 116.200 ;
        RECT 175.800 115.800 202.600 116.100 ;
        RECT 11.000 114.800 11.400 115.200 ;
        RECT 20.600 115.100 21.000 115.200 ;
        RECT 22.200 115.100 22.500 115.800 ;
        RECT 20.600 114.800 22.500 115.100 ;
        RECT 27.000 114.800 27.400 115.200 ;
        RECT 30.200 115.100 30.600 115.200 ;
        RECT 38.200 115.100 38.600 115.200 ;
        RECT 30.200 114.800 38.600 115.100 ;
        RECT 41.400 115.100 41.800 115.200 ;
        RECT 42.200 115.100 42.600 115.200 ;
        RECT 41.400 114.800 42.600 115.100 ;
        RECT 43.800 115.100 44.200 115.200 ;
        RECT 76.600 115.100 77.000 115.200 ;
        RECT 79.800 115.100 80.200 115.200 ;
        RECT 43.800 114.800 64.900 115.100 ;
        RECT 76.600 114.800 80.200 115.100 ;
        RECT 86.200 115.100 86.600 115.200 ;
        RECT 95.800 115.100 96.200 115.200 ;
        RECT 99.800 115.100 100.200 115.200 ;
        RECT 86.200 114.800 100.200 115.100 ;
        RECT 105.400 115.100 105.800 115.200 ;
        RECT 109.400 115.100 109.700 115.800 ;
        RECT 138.200 115.200 138.500 115.800 ;
        RECT 105.400 114.800 109.700 115.100 ;
        RECT 129.400 115.100 129.800 115.200 ;
        RECT 130.200 115.100 130.600 115.200 ;
        RECT 129.400 114.800 130.600 115.100 ;
        RECT 138.200 114.800 138.600 115.200 ;
        RECT 143.800 114.800 144.200 115.200 ;
        RECT 151.000 115.100 151.400 115.200 ;
        RECT 156.600 115.100 157.000 115.200 ;
        RECT 160.600 115.100 161.000 115.200 ;
        RECT 151.000 114.800 161.000 115.100 ;
        RECT 164.600 114.800 165.000 115.200 ;
        RECT 199.000 115.100 199.400 115.200 ;
        RECT 191.000 114.800 199.400 115.100 ;
        RECT 3.000 114.100 3.400 114.200 ;
        RECT 11.000 114.100 11.300 114.800 ;
        RECT 27.000 114.100 27.300 114.800 ;
        RECT 3.000 113.800 27.300 114.100 ;
        RECT 42.200 114.100 42.600 114.200 ;
        RECT 47.000 114.100 47.400 114.200 ;
        RECT 42.200 113.800 47.400 114.100 ;
        RECT 48.600 114.100 49.000 114.200 ;
        RECT 51.800 114.100 52.200 114.200 ;
        RECT 54.200 114.100 54.600 114.200 ;
        RECT 55.800 114.100 56.200 114.200 ;
        RECT 48.600 113.800 56.200 114.100 ;
        RECT 60.600 114.100 61.000 114.200 ;
        RECT 63.800 114.100 64.200 114.200 ;
        RECT 60.600 113.800 64.200 114.100 ;
        RECT 64.600 114.100 64.900 114.800 ;
        RECT 89.400 114.100 89.800 114.200 ;
        RECT 64.600 113.800 89.800 114.100 ;
        RECT 105.400 114.100 105.800 114.200 ;
        RECT 107.800 114.100 108.200 114.200 ;
        RECT 111.000 114.100 111.400 114.200 ;
        RECT 105.400 113.800 111.400 114.100 ;
        RECT 117.400 114.100 117.800 114.200 ;
        RECT 118.200 114.100 118.600 114.200 ;
        RECT 117.400 113.800 118.600 114.100 ;
        RECT 125.400 114.100 125.800 114.200 ;
        RECT 129.400 114.100 129.800 114.200 ;
        RECT 125.400 113.800 129.800 114.100 ;
        RECT 131.000 114.100 131.400 114.200 ;
        RECT 131.800 114.100 132.200 114.200 ;
        RECT 131.000 113.800 132.200 114.100 ;
        RECT 143.800 114.100 144.100 114.800 ;
        RECT 164.600 114.200 164.900 114.800 ;
        RECT 191.000 114.200 191.300 114.800 ;
        RECT 157.400 114.100 157.800 114.200 ;
        RECT 160.600 114.100 161.000 114.200 ;
        RECT 162.200 114.100 162.600 114.200 ;
        RECT 143.800 113.800 156.900 114.100 ;
        RECT 157.400 113.800 162.600 114.100 ;
        RECT 164.600 113.800 165.000 114.200 ;
        RECT 175.800 114.100 176.200 114.200 ;
        RECT 188.600 114.100 189.000 114.200 ;
        RECT 175.800 113.800 189.000 114.100 ;
        RECT 191.000 113.800 191.400 114.200 ;
        RECT 14.200 113.100 14.600 113.200 ;
        RECT 23.000 113.100 23.400 113.200 ;
        RECT 14.200 112.800 23.400 113.100 ;
        RECT 37.400 113.100 37.800 113.200 ;
        RECT 40.600 113.100 41.000 113.200 ;
        RECT 47.800 113.100 48.200 113.200 ;
        RECT 37.400 112.800 48.200 113.100 ;
        RECT 52.600 113.100 53.000 113.200 ;
        RECT 61.400 113.100 61.800 113.200 ;
        RECT 52.600 112.800 61.800 113.100 ;
        RECT 63.800 113.100 64.200 113.200 ;
        RECT 67.800 113.100 68.200 113.200 ;
        RECT 76.600 113.100 77.000 113.200 ;
        RECT 63.800 112.800 77.000 113.100 ;
        RECT 97.400 113.100 97.800 113.200 ;
        RECT 102.200 113.100 102.600 113.200 ;
        RECT 97.400 112.800 102.600 113.100 ;
        RECT 115.800 113.100 116.200 113.200 ;
        RECT 126.200 113.100 126.600 113.200 ;
        RECT 115.800 112.800 126.600 113.100 ;
        RECT 131.000 113.100 131.400 113.200 ;
        RECT 146.200 113.100 146.600 113.200 ;
        RECT 131.000 112.800 146.600 113.100 ;
        RECT 155.800 112.800 156.200 113.200 ;
        RECT 156.600 113.100 156.900 113.800 ;
        RECT 163.800 113.100 164.200 113.200 ;
        RECT 165.400 113.100 165.800 113.200 ;
        RECT 156.600 112.800 159.300 113.100 ;
        RECT 163.800 112.800 165.800 113.100 ;
        RECT 175.000 113.100 175.400 113.200 ;
        RECT 175.800 113.100 176.100 113.800 ;
        RECT 175.000 112.800 176.100 113.100 ;
        RECT 61.400 112.100 61.700 112.800 ;
        RECT 65.400 112.100 65.800 112.200 ;
        RECT 67.800 112.100 68.200 112.200 ;
        RECT 61.400 111.800 68.200 112.100 ;
        RECT 82.200 112.100 82.600 112.200 ;
        RECT 112.600 112.100 113.000 112.200 ;
        RECT 82.200 111.800 113.000 112.100 ;
        RECT 115.000 112.100 115.400 112.200 ;
        RECT 120.600 112.100 121.000 112.200 ;
        RECT 133.400 112.100 133.800 112.200 ;
        RECT 115.000 111.800 133.800 112.100 ;
        RECT 155.800 112.100 156.100 112.800 ;
        RECT 159.000 112.200 159.300 112.800 ;
        RECT 158.200 112.100 158.600 112.200 ;
        RECT 155.800 111.800 158.600 112.100 ;
        RECT 159.000 111.800 159.400 112.200 ;
        RECT 163.800 112.100 164.200 112.200 ;
        RECT 194.200 112.100 194.600 112.200 ;
        RECT 198.200 112.100 198.600 112.200 ;
        RECT 163.800 111.800 198.600 112.100 ;
        RECT 45.400 111.100 45.800 111.200 ;
        RECT 48.600 111.100 49.000 111.200 ;
        RECT 45.400 110.800 49.000 111.100 ;
        RECT 55.000 111.100 55.400 111.200 ;
        RECT 70.200 111.100 70.600 111.200 ;
        RECT 55.000 110.800 70.600 111.100 ;
        RECT 124.600 111.100 125.000 111.200 ;
        RECT 127.000 111.100 127.400 111.200 ;
        RECT 124.600 110.800 127.400 111.100 ;
        RECT 128.600 111.100 129.000 111.200 ;
        RECT 196.600 111.100 197.000 111.200 ;
        RECT 128.600 110.800 197.000 111.100 ;
        RECT 16.600 110.100 17.000 110.200 ;
        RECT 39.800 110.100 40.200 110.200 ;
        RECT 16.600 109.800 40.200 110.100 ;
        RECT 47.000 110.100 47.400 110.200 ;
        RECT 55.000 110.100 55.400 110.200 ;
        RECT 58.200 110.100 58.600 110.200 ;
        RECT 47.000 109.800 58.600 110.100 ;
        RECT 64.600 110.100 65.000 110.200 ;
        RECT 67.000 110.100 67.400 110.200 ;
        RECT 64.600 109.800 67.400 110.100 ;
        RECT 71.000 110.100 71.400 110.200 ;
        RECT 71.800 110.100 72.200 110.200 ;
        RECT 71.000 109.800 72.200 110.100 ;
        RECT 72.600 110.100 73.000 110.200 ;
        RECT 82.200 110.100 82.600 110.200 ;
        RECT 72.600 109.800 82.600 110.100 ;
        RECT 123.800 110.100 124.200 110.200 ;
        RECT 127.800 110.100 128.200 110.200 ;
        RECT 151.000 110.100 151.400 110.200 ;
        RECT 123.800 109.800 151.400 110.100 ;
        RECT 155.800 110.100 156.200 110.200 ;
        RECT 162.200 110.100 162.600 110.200 ;
        RECT 155.800 109.800 162.600 110.100 ;
        RECT 185.400 110.100 185.800 110.200 ;
        RECT 193.400 110.100 193.800 110.200 ;
        RECT 201.400 110.100 201.800 110.200 ;
        RECT 185.400 109.800 201.800 110.100 ;
        RECT 5.400 109.100 5.800 109.200 ;
        RECT 18.200 109.100 18.600 109.200 ;
        RECT 5.400 108.800 18.600 109.100 ;
        RECT 22.200 108.800 22.600 109.200 ;
        RECT 35.800 109.100 36.200 109.200 ;
        RECT 27.800 108.800 36.200 109.100 ;
        RECT 41.400 109.100 41.800 109.200 ;
        RECT 57.400 109.100 57.800 109.200 ;
        RECT 41.400 108.800 57.800 109.100 ;
        RECT 64.600 108.800 65.000 109.200 ;
        RECT 70.200 109.100 70.600 109.200 ;
        RECT 83.000 109.100 83.400 109.200 ;
        RECT 70.200 108.800 83.400 109.100 ;
        RECT 85.400 109.100 85.800 109.200 ;
        RECT 87.800 109.100 88.200 109.200 ;
        RECT 90.200 109.100 90.600 109.200 ;
        RECT 85.400 108.800 90.600 109.100 ;
        RECT 94.200 108.800 94.600 109.200 ;
        RECT 121.400 109.100 121.800 109.200 ;
        RECT 131.800 109.100 132.200 109.200 ;
        RECT 121.400 108.800 132.200 109.100 ;
        RECT 159.800 108.800 160.200 109.200 ;
        RECT 167.800 108.800 168.200 109.200 ;
        RECT 171.000 108.800 171.400 109.200 ;
        RECT 172.600 109.100 173.000 109.200 ;
        RECT 173.400 109.100 173.800 109.200 ;
        RECT 172.600 108.800 173.800 109.100 ;
        RECT 0.600 108.100 1.000 108.200 ;
        RECT 17.400 108.100 17.800 108.200 ;
        RECT 22.200 108.100 22.500 108.800 ;
        RECT 27.800 108.200 28.100 108.800 ;
        RECT 64.600 108.200 64.900 108.800 ;
        RECT 0.600 107.800 22.500 108.100 ;
        RECT 25.400 108.100 25.800 108.200 ;
        RECT 26.200 108.100 26.600 108.200 ;
        RECT 25.400 107.800 26.600 108.100 ;
        RECT 27.800 107.800 28.200 108.200 ;
        RECT 31.000 108.100 31.400 108.200 ;
        RECT 31.800 108.100 32.200 108.200 ;
        RECT 31.000 107.800 32.200 108.100 ;
        RECT 39.800 108.100 40.200 108.200 ;
        RECT 40.600 108.100 41.000 108.200 ;
        RECT 39.800 107.800 41.000 108.100 ;
        RECT 41.400 108.100 41.800 108.200 ;
        RECT 43.800 108.100 44.200 108.200 ;
        RECT 41.400 107.800 44.200 108.100 ;
        RECT 46.200 108.100 46.600 108.200 ;
        RECT 47.000 108.100 47.400 108.200 ;
        RECT 46.200 107.800 47.400 108.100 ;
        RECT 64.600 107.800 65.000 108.200 ;
        RECT 68.600 108.100 69.000 108.200 ;
        RECT 69.400 108.100 69.800 108.200 ;
        RECT 68.600 107.800 69.800 108.100 ;
        RECT 71.800 108.100 72.200 108.200 ;
        RECT 72.600 108.100 73.000 108.200 ;
        RECT 71.800 107.800 73.000 108.100 ;
        RECT 79.800 108.100 80.200 108.200 ;
        RECT 88.600 108.100 89.000 108.200 ;
        RECT 79.800 107.800 89.000 108.100 ;
        RECT 90.200 108.100 90.600 108.200 ;
        RECT 94.200 108.100 94.500 108.800 ;
        RECT 90.200 107.800 94.500 108.100 ;
        RECT 113.400 107.800 113.800 108.200 ;
        RECT 129.400 108.100 129.800 108.200 ;
        RECT 134.200 108.100 134.600 108.200 ;
        RECT 137.400 108.100 137.800 108.200 ;
        RECT 129.400 107.800 137.800 108.100 ;
        RECT 159.800 108.100 160.100 108.800 ;
        RECT 164.600 108.100 165.000 108.200 ;
        RECT 159.800 107.800 165.000 108.100 ;
        RECT 166.200 108.100 166.600 108.200 ;
        RECT 167.800 108.100 168.100 108.800 ;
        RECT 166.200 107.800 168.100 108.100 ;
        RECT 169.400 108.100 169.800 108.200 ;
        RECT 170.200 108.100 170.600 108.200 ;
        RECT 169.400 107.800 170.600 108.100 ;
        RECT 171.000 108.100 171.300 108.800 ;
        RECT 175.000 108.100 175.400 108.200 ;
        RECT 171.000 107.800 175.400 108.100 ;
        RECT 176.600 108.100 177.000 108.200 ;
        RECT 192.600 108.100 193.000 108.200 ;
        RECT 176.600 107.800 193.000 108.100 ;
        RECT 12.600 107.100 13.000 107.200 ;
        RECT 17.400 107.100 17.800 107.200 ;
        RECT 12.600 106.800 17.800 107.100 ;
        RECT 24.600 107.100 25.000 107.200 ;
        RECT 30.200 107.100 30.600 107.200 ;
        RECT 35.000 107.100 35.400 107.200 ;
        RECT 37.400 107.100 37.800 107.200 ;
        RECT 42.200 107.100 42.600 107.200 ;
        RECT 45.400 107.100 45.800 107.200 ;
        RECT 24.600 106.800 45.800 107.100 ;
        RECT 51.000 107.100 51.400 107.200 ;
        RECT 54.200 107.100 54.600 107.200 ;
        RECT 51.000 106.800 54.600 107.100 ;
        RECT 57.400 106.800 57.800 107.200 ;
        RECT 67.000 107.100 67.400 107.200 ;
        RECT 75.000 107.100 75.400 107.200 ;
        RECT 89.400 107.100 89.800 107.200 ;
        RECT 67.000 106.800 75.400 107.100 ;
        RECT 87.000 106.800 89.800 107.100 ;
        RECT 92.600 107.100 93.000 107.200 ;
        RECT 93.400 107.100 93.800 107.200 ;
        RECT 92.600 106.800 93.800 107.100 ;
        RECT 99.800 107.100 100.200 107.200 ;
        RECT 104.600 107.100 105.000 107.200 ;
        RECT 99.800 106.800 105.000 107.100 ;
        RECT 113.400 107.100 113.700 107.800 ;
        RECT 120.600 107.100 121.000 107.200 ;
        RECT 113.400 106.800 121.000 107.100 ;
        RECT 129.400 107.100 129.800 107.200 ;
        RECT 132.600 107.100 133.000 107.200 ;
        RECT 135.800 107.100 136.200 107.200 ;
        RECT 129.400 106.800 136.200 107.100 ;
        RECT 136.600 107.100 137.000 107.200 ;
        RECT 145.400 107.100 145.800 107.200 ;
        RECT 136.600 106.800 145.800 107.100 ;
        RECT 147.000 107.100 147.400 107.200 ;
        RECT 160.600 107.100 161.000 107.200 ;
        RECT 163.800 107.100 164.200 107.200 ;
        RECT 147.000 106.800 164.200 107.100 ;
        RECT 165.400 107.100 165.800 107.200 ;
        RECT 187.000 107.100 187.400 107.200 ;
        RECT 165.400 106.800 187.400 107.100 ;
        RECT 197.400 107.100 197.800 107.200 ;
        RECT 199.800 107.100 200.200 107.200 ;
        RECT 197.400 106.800 200.200 107.100 ;
        RECT 57.400 106.200 57.700 106.800 ;
        RECT 87.000 106.200 87.300 106.800 ;
        RECT 13.400 106.100 13.800 106.200 ;
        RECT 15.000 106.100 15.400 106.200 ;
        RECT 13.400 105.800 15.400 106.100 ;
        RECT 27.000 106.100 27.400 106.200 ;
        RECT 32.600 106.100 33.000 106.200 ;
        RECT 41.400 106.100 41.800 106.200 ;
        RECT 27.000 105.800 32.100 106.100 ;
        RECT 32.600 105.800 41.800 106.100 ;
        RECT 42.200 105.800 42.600 106.200 ;
        RECT 43.000 105.800 43.400 106.200 ;
        RECT 51.800 106.100 52.200 106.200 ;
        RECT 52.600 106.100 53.000 106.200 ;
        RECT 51.800 105.800 53.000 106.100 ;
        RECT 57.400 105.800 57.800 106.200 ;
        RECT 68.600 106.100 69.000 106.200 ;
        RECT 69.400 106.100 69.800 106.200 ;
        RECT 68.600 105.800 69.800 106.100 ;
        RECT 72.600 106.100 73.000 106.200 ;
        RECT 85.400 106.100 85.800 106.200 ;
        RECT 72.600 105.800 85.800 106.100 ;
        RECT 87.000 105.800 87.400 106.200 ;
        RECT 95.800 106.100 96.200 106.200 ;
        RECT 96.600 106.100 97.000 106.200 ;
        RECT 102.200 106.100 102.600 106.200 ;
        RECT 110.200 106.100 110.600 106.200 ;
        RECT 95.800 105.800 102.600 106.100 ;
        RECT 103.000 105.800 110.600 106.100 ;
        RECT 123.800 106.100 124.200 106.200 ;
        RECT 137.400 106.100 137.800 106.200 ;
        RECT 160.600 106.100 161.000 106.200 ;
        RECT 123.800 105.800 133.700 106.100 ;
        RECT 137.400 105.800 161.000 106.100 ;
        RECT 165.400 106.100 165.800 106.200 ;
        RECT 170.200 106.100 170.600 106.200 ;
        RECT 171.000 106.100 171.400 106.200 ;
        RECT 165.400 105.800 171.400 106.100 ;
        RECT 171.800 106.100 172.200 106.200 ;
        RECT 172.600 106.100 173.000 106.200 ;
        RECT 171.800 105.800 173.000 106.100 ;
        RECT 191.000 106.100 191.400 106.200 ;
        RECT 192.600 106.100 193.000 106.200 ;
        RECT 195.000 106.100 195.400 106.200 ;
        RECT 191.000 105.800 195.400 106.100 ;
        RECT 31.800 105.200 32.100 105.800 ;
        RECT 42.200 105.200 42.500 105.800 ;
        RECT 43.000 105.200 43.300 105.800 ;
        RECT 103.000 105.200 103.300 105.800 ;
        RECT 133.400 105.200 133.700 105.800 ;
        RECT 7.000 105.100 7.400 105.200 ;
        RECT 7.000 104.800 12.900 105.100 ;
        RECT 12.600 104.200 12.900 104.800 ;
        RECT 21.400 104.800 21.800 105.200 ;
        RECT 31.800 104.800 32.200 105.200 ;
        RECT 42.200 104.800 42.600 105.200 ;
        RECT 43.000 104.800 43.400 105.200 ;
        RECT 67.800 105.100 68.200 105.200 ;
        RECT 69.400 105.100 69.800 105.200 ;
        RECT 67.800 104.800 69.800 105.100 ;
        RECT 85.400 104.800 85.800 105.200 ;
        RECT 91.000 105.100 91.400 105.200 ;
        RECT 97.400 105.100 97.800 105.200 ;
        RECT 91.000 104.800 97.800 105.100 ;
        RECT 103.000 104.800 103.400 105.200 ;
        RECT 133.400 105.100 133.800 105.200 ;
        RECT 135.000 105.100 135.400 105.200 ;
        RECT 133.400 104.800 135.400 105.100 ;
        RECT 179.800 105.100 180.200 105.200 ;
        RECT 180.600 105.100 181.000 105.200 ;
        RECT 179.800 104.800 181.000 105.100 ;
        RECT 183.800 105.100 184.200 105.200 ;
        RECT 195.000 105.100 195.400 105.200 ;
        RECT 183.800 104.800 195.400 105.100 ;
        RECT 21.400 104.200 21.700 104.800 ;
        RECT 85.400 104.200 85.700 104.800 ;
        RECT 11.000 103.800 11.400 104.200 ;
        RECT 12.600 103.800 13.000 104.200 ;
        RECT 21.400 103.800 21.800 104.200 ;
        RECT 27.000 104.100 27.400 104.200 ;
        RECT 33.400 104.100 33.800 104.200 ;
        RECT 27.000 103.800 33.800 104.100 ;
        RECT 39.800 104.100 40.200 104.200 ;
        RECT 43.800 104.100 44.200 104.200 ;
        RECT 39.800 103.800 44.200 104.100 ;
        RECT 56.600 104.100 57.000 104.200 ;
        RECT 69.400 104.100 69.800 104.200 ;
        RECT 56.600 103.800 69.800 104.100 ;
        RECT 85.400 103.800 85.800 104.200 ;
        RECT 90.200 104.100 90.600 104.200 ;
        RECT 91.800 104.100 92.200 104.200 ;
        RECT 90.200 103.800 92.200 104.100 ;
        RECT 98.200 104.100 98.600 104.200 ;
        RECT 104.600 104.100 105.000 104.200 ;
        RECT 98.200 103.800 105.000 104.100 ;
        RECT 112.600 104.100 113.000 104.200 ;
        RECT 121.400 104.100 121.800 104.200 ;
        RECT 139.800 104.100 140.200 104.200 ;
        RECT 112.600 103.800 140.200 104.100 ;
        RECT 182.200 104.100 182.600 104.200 ;
        RECT 187.800 104.100 188.200 104.200 ;
        RECT 182.200 103.800 188.200 104.100 ;
        RECT 11.000 103.100 11.300 103.800 ;
        RECT 20.600 103.100 21.000 103.200 ;
        RECT 37.400 103.100 37.800 103.200 ;
        RECT 11.000 102.800 37.800 103.100 ;
        RECT 55.800 103.100 56.200 103.200 ;
        RECT 91.000 103.100 91.400 103.200 ;
        RECT 55.800 102.800 91.400 103.100 ;
        RECT 113.400 103.100 113.800 103.200 ;
        RECT 114.200 103.100 114.600 103.200 ;
        RECT 113.400 102.800 114.600 103.100 ;
        RECT 116.600 103.100 117.000 103.200 ;
        RECT 117.400 103.100 117.800 103.200 ;
        RECT 154.200 103.100 154.600 103.200 ;
        RECT 116.600 102.800 154.600 103.100 ;
        RECT 160.600 103.100 161.000 103.200 ;
        RECT 190.200 103.100 190.600 103.200 ;
        RECT 160.600 102.800 190.600 103.100 ;
        RECT 200.600 103.100 201.000 103.200 ;
        RECT 202.200 103.100 202.600 103.200 ;
        RECT 200.600 102.800 202.600 103.100 ;
        RECT 58.200 102.100 58.600 102.200 ;
        RECT 73.400 102.100 73.800 102.200 ;
        RECT 58.200 101.800 73.800 102.100 ;
        RECT 80.600 101.800 81.000 102.200 ;
        RECT 132.600 102.100 133.000 102.200 ;
        RECT 136.600 102.100 137.000 102.200 ;
        RECT 132.600 101.800 137.000 102.100 ;
        RECT 148.600 102.100 149.000 102.200 ;
        RECT 202.200 102.100 202.600 102.200 ;
        RECT 148.600 101.800 202.600 102.100 ;
        RECT 80.600 101.200 80.900 101.800 ;
        RECT 60.600 101.100 61.000 101.200 ;
        RECT 75.800 101.100 76.200 101.200 ;
        RECT 60.600 100.800 76.200 101.100 ;
        RECT 80.600 101.100 81.000 101.200 ;
        RECT 89.400 101.100 89.800 101.200 ;
        RECT 80.600 100.800 89.800 101.100 ;
        RECT 102.200 101.100 102.600 101.200 ;
        RECT 126.200 101.100 126.600 101.200 ;
        RECT 102.200 100.800 126.600 101.100 ;
        RECT 190.200 101.100 190.600 101.200 ;
        RECT 191.000 101.100 191.400 101.200 ;
        RECT 190.200 100.800 191.400 101.100 ;
        RECT 62.200 99.800 62.600 100.200 ;
        RECT 64.600 100.100 65.000 100.200 ;
        RECT 71.800 100.100 72.200 100.200 ;
        RECT 76.600 100.100 77.000 100.200 ;
        RECT 127.800 100.100 128.200 100.200 ;
        RECT 64.600 99.800 77.000 100.100 ;
        RECT 115.800 99.800 128.200 100.100 ;
        RECT 169.400 99.800 169.800 100.200 ;
        RECT 62.200 99.200 62.500 99.800 ;
        RECT 27.800 99.100 28.200 99.200 ;
        RECT 38.200 99.100 38.600 99.200 ;
        RECT 27.800 98.800 38.600 99.100 ;
        RECT 40.600 99.100 41.000 99.200 ;
        RECT 47.800 99.100 48.200 99.200 ;
        RECT 40.600 98.800 48.200 99.100 ;
        RECT 62.200 98.800 62.600 99.200 ;
        RECT 71.800 99.100 72.200 99.200 ;
        RECT 78.200 99.100 78.600 99.200 ;
        RECT 71.800 98.800 78.600 99.100 ;
        RECT 81.400 98.800 81.800 99.200 ;
        RECT 87.000 99.100 87.400 99.200 ;
        RECT 93.400 99.100 93.800 99.200 ;
        RECT 115.800 99.100 116.100 99.800 ;
        RECT 169.400 99.200 169.700 99.800 ;
        RECT 87.000 98.800 116.100 99.100 ;
        RECT 123.800 99.100 124.200 99.200 ;
        RECT 125.400 99.100 125.800 99.200 ;
        RECT 144.600 99.100 145.000 99.200 ;
        RECT 148.600 99.100 149.000 99.200 ;
        RECT 150.200 99.100 150.600 99.200 ;
        RECT 123.800 98.800 150.600 99.100 ;
        RECT 169.400 98.800 169.800 99.200 ;
        RECT 47.800 98.100 48.200 98.200 ;
        RECT 30.200 97.800 48.200 98.100 ;
        RECT 74.200 97.800 74.600 98.200 ;
        RECT 75.800 98.100 76.200 98.200 ;
        RECT 81.400 98.100 81.700 98.800 ;
        RECT 75.800 97.800 81.700 98.100 ;
        RECT 86.200 97.800 86.600 98.200 ;
        RECT 91.800 98.100 92.200 98.200 ;
        RECT 92.600 98.100 93.000 98.200 ;
        RECT 91.800 97.800 93.000 98.100 ;
        RECT 99.000 98.100 99.400 98.200 ;
        RECT 115.000 98.100 115.400 98.200 ;
        RECT 99.000 97.800 115.400 98.100 ;
        RECT 116.600 98.100 117.000 98.200 ;
        RECT 123.800 98.100 124.100 98.800 ;
        RECT 116.600 97.800 124.100 98.100 ;
        RECT 151.800 98.100 152.200 98.200 ;
        RECT 167.800 98.100 168.200 98.200 ;
        RECT 151.800 97.800 168.200 98.100 ;
        RECT 30.200 97.200 30.500 97.800 ;
        RECT 74.200 97.200 74.500 97.800 ;
        RECT 86.200 97.200 86.500 97.800 ;
        RECT 30.200 96.800 30.600 97.200 ;
        RECT 36.600 96.800 37.000 97.200 ;
        RECT 49.400 97.100 49.800 97.200 ;
        RECT 53.400 97.100 53.800 97.200 ;
        RECT 58.200 97.100 58.600 97.200 ;
        RECT 49.400 96.800 58.600 97.100 ;
        RECT 65.400 97.100 65.800 97.200 ;
        RECT 72.600 97.100 73.000 97.200 ;
        RECT 65.400 96.800 73.000 97.100 ;
        RECT 74.200 96.800 74.600 97.200 ;
        RECT 76.600 97.100 77.000 97.200 ;
        RECT 79.000 97.100 79.400 97.200 ;
        RECT 83.000 97.100 83.400 97.200 ;
        RECT 76.600 96.800 83.400 97.100 ;
        RECT 86.200 96.800 86.600 97.200 ;
        RECT 107.800 97.100 108.200 97.200 ;
        RECT 118.200 97.100 118.600 97.200 ;
        RECT 107.800 96.800 118.600 97.100 ;
        RECT 126.200 97.100 126.600 97.200 ;
        RECT 161.400 97.100 161.800 97.200 ;
        RECT 126.200 96.800 161.800 97.100 ;
        RECT 162.200 97.100 162.600 97.200 ;
        RECT 162.200 96.800 172.100 97.100 ;
        RECT 18.200 96.100 18.600 96.200 ;
        RECT 22.200 96.100 22.600 96.200 ;
        RECT 23.000 96.100 23.400 96.200 ;
        RECT 18.200 95.800 23.400 96.100 ;
        RECT 36.600 96.100 36.900 96.800 ;
        RECT 171.800 96.200 172.100 96.800 ;
        RECT 39.800 96.100 40.200 96.200 ;
        RECT 36.600 95.800 40.200 96.100 ;
        RECT 41.400 96.100 41.800 96.200 ;
        RECT 45.400 96.100 45.800 96.200 ;
        RECT 41.400 95.800 45.800 96.100 ;
        RECT 47.000 96.100 47.400 96.200 ;
        RECT 119.800 96.100 120.200 96.200 ;
        RECT 122.200 96.100 122.600 96.200 ;
        RECT 163.000 96.100 163.400 96.200 ;
        RECT 166.200 96.100 166.600 96.200 ;
        RECT 47.000 95.800 166.600 96.100 ;
        RECT 169.400 95.800 169.800 96.200 ;
        RECT 171.800 95.800 172.200 96.200 ;
        RECT 180.600 96.100 181.000 96.200 ;
        RECT 200.600 96.100 201.000 96.200 ;
        RECT 179.800 95.800 201.000 96.100 ;
        RECT 12.600 95.100 13.000 95.200 ;
        RECT 19.800 95.100 20.200 95.200 ;
        RECT 12.600 94.800 20.200 95.100 ;
        RECT 20.600 94.800 21.000 95.200 ;
        RECT 31.800 94.800 32.200 95.200 ;
        RECT 33.400 95.100 33.800 95.200 ;
        RECT 55.000 95.100 55.400 95.200 ;
        RECT 64.600 95.100 65.000 95.200 ;
        RECT 66.200 95.100 66.600 95.200 ;
        RECT 33.400 94.800 54.500 95.100 ;
        RECT 55.000 94.800 66.600 95.100 ;
        RECT 73.400 95.100 73.800 95.200 ;
        RECT 79.000 95.100 79.400 95.200 ;
        RECT 83.000 95.100 83.400 95.200 ;
        RECT 73.400 94.800 74.500 95.100 ;
        RECT 79.000 94.800 83.400 95.100 ;
        RECT 85.400 95.100 85.800 95.200 ;
        RECT 93.400 95.100 93.800 95.200 ;
        RECT 96.600 95.100 97.000 95.200 ;
        RECT 85.400 94.800 97.000 95.100 ;
        RECT 105.400 95.100 105.800 95.200 ;
        RECT 108.600 95.100 109.000 95.200 ;
        RECT 105.400 94.800 109.000 95.100 ;
        RECT 113.400 95.100 113.800 95.200 ;
        RECT 115.800 95.100 116.200 95.200 ;
        RECT 117.400 95.100 117.800 95.200 ;
        RECT 113.400 94.800 117.800 95.100 ;
        RECT 138.200 95.100 138.600 95.200 ;
        RECT 139.000 95.100 139.400 95.200 ;
        RECT 138.200 94.800 139.400 95.100 ;
        RECT 139.800 95.100 140.200 95.200 ;
        RECT 141.400 95.100 141.800 95.200 ;
        RECT 139.800 94.800 141.800 95.100 ;
        RECT 145.400 94.800 145.800 95.200 ;
        RECT 146.200 95.100 146.600 95.200 ;
        RECT 156.600 95.100 157.000 95.200 ;
        RECT 167.000 95.100 167.400 95.200 ;
        RECT 146.200 94.800 167.400 95.100 ;
        RECT 169.400 95.100 169.700 95.800 ;
        RECT 182.200 95.100 182.600 95.200 ;
        RECT 169.400 94.800 182.600 95.100 ;
        RECT 15.800 94.100 16.200 94.200 ;
        RECT 20.600 94.100 20.900 94.800 ;
        RECT 31.800 94.100 32.100 94.800 ;
        RECT 15.800 93.800 32.100 94.100 ;
        RECT 33.400 93.800 33.800 94.200 ;
        RECT 45.400 94.100 45.800 94.200 ;
        RECT 46.200 94.100 46.600 94.200 ;
        RECT 45.400 93.800 46.600 94.100 ;
        RECT 47.800 94.100 48.200 94.200 ;
        RECT 48.600 94.100 49.000 94.200 ;
        RECT 47.800 93.800 49.000 94.100 ;
        RECT 53.400 93.800 53.800 94.200 ;
        RECT 54.200 94.100 54.500 94.800 ;
        RECT 74.200 94.200 74.500 94.800 ;
        RECT 145.400 94.200 145.700 94.800 ;
        RECT 57.400 94.100 57.800 94.200 ;
        RECT 54.200 93.800 57.800 94.100 ;
        RECT 59.000 94.100 59.400 94.200 ;
        RECT 59.800 94.100 60.200 94.200 ;
        RECT 59.000 93.800 60.200 94.100 ;
        RECT 63.800 94.100 64.200 94.200 ;
        RECT 64.600 94.100 65.000 94.200 ;
        RECT 63.800 93.800 65.000 94.100 ;
        RECT 74.200 93.800 74.600 94.200 ;
        RECT 78.200 94.100 78.600 94.200 ;
        RECT 79.800 94.100 80.200 94.200 ;
        RECT 78.200 93.800 80.200 94.100 ;
        RECT 82.200 94.100 82.600 94.200 ;
        RECT 99.000 94.100 99.400 94.200 ;
        RECT 82.200 93.800 99.400 94.100 ;
        RECT 99.800 94.100 100.200 94.200 ;
        RECT 112.600 94.100 113.000 94.200 ;
        RECT 123.000 94.100 123.400 94.200 ;
        RECT 99.800 93.800 123.400 94.100 ;
        RECT 127.000 94.100 127.400 94.200 ;
        RECT 138.200 94.100 138.600 94.200 ;
        RECT 143.800 94.100 144.200 94.200 ;
        RECT 127.000 93.800 130.500 94.100 ;
        RECT 138.200 93.800 144.200 94.100 ;
        RECT 145.400 93.800 145.800 94.200 ;
        RECT 147.000 94.100 147.400 94.200 ;
        RECT 149.400 94.100 149.800 94.200 ;
        RECT 147.000 93.800 149.800 94.100 ;
        RECT 150.200 94.100 150.600 94.200 ;
        RECT 151.000 94.100 151.400 94.200 ;
        RECT 150.200 93.800 151.400 94.100 ;
        RECT 152.600 93.800 153.000 94.200 ;
        RECT 162.200 94.100 162.600 94.200 ;
        RECT 160.600 93.800 162.600 94.100 ;
        RECT 165.400 94.100 165.800 94.200 ;
        RECT 166.200 94.100 166.600 94.200 ;
        RECT 165.400 93.800 166.600 94.100 ;
        RECT 171.000 94.100 171.400 94.200 ;
        RECT 175.000 94.100 175.400 94.200 ;
        RECT 171.000 93.800 175.400 94.100 ;
        RECT 189.400 94.100 189.800 94.200 ;
        RECT 198.200 94.100 198.600 94.200 ;
        RECT 189.400 93.800 198.600 94.100 ;
        RECT 27.000 93.100 27.400 93.200 ;
        RECT 28.600 93.100 29.000 93.200 ;
        RECT 27.000 92.800 29.000 93.100 ;
        RECT 33.400 93.100 33.700 93.800 ;
        RECT 35.800 93.100 36.200 93.200 ;
        RECT 33.400 92.800 36.200 93.100 ;
        RECT 39.800 93.100 40.200 93.200 ;
        RECT 40.600 93.100 41.000 93.200 ;
        RECT 39.800 92.800 41.000 93.100 ;
        RECT 42.200 93.100 42.600 93.200 ;
        RECT 53.400 93.100 53.700 93.800 ;
        RECT 130.200 93.200 130.500 93.800 ;
        RECT 42.200 92.800 53.700 93.100 ;
        RECT 75.800 93.100 76.200 93.200 ;
        RECT 83.800 93.100 84.200 93.200 ;
        RECT 75.800 92.800 84.200 93.100 ;
        RECT 84.600 93.100 85.000 93.200 ;
        RECT 85.400 93.100 85.800 93.200 ;
        RECT 84.600 92.800 85.800 93.100 ;
        RECT 89.400 93.100 89.800 93.200 ;
        RECT 90.200 93.100 90.600 93.200 ;
        RECT 89.400 92.800 90.600 93.100 ;
        RECT 91.000 93.100 91.400 93.200 ;
        RECT 115.800 93.100 116.200 93.200 ;
        RECT 91.000 92.800 116.200 93.100 ;
        RECT 130.200 92.800 130.600 93.200 ;
        RECT 132.600 93.100 133.000 93.200 ;
        RECT 143.800 93.100 144.200 93.200 ;
        RECT 147.800 93.100 148.200 93.200 ;
        RECT 132.600 92.800 140.900 93.100 ;
        RECT 143.800 92.800 148.200 93.100 ;
        RECT 151.000 93.100 151.400 93.200 ;
        RECT 152.600 93.100 152.900 93.800 ;
        RECT 160.600 93.200 160.900 93.800 ;
        RECT 151.000 92.800 152.900 93.100 ;
        RECT 154.200 93.100 154.600 93.200 ;
        RECT 155.000 93.100 155.400 93.200 ;
        RECT 154.200 92.800 155.400 93.100 ;
        RECT 159.000 93.100 159.400 93.200 ;
        RECT 159.800 93.100 160.200 93.200 ;
        RECT 159.000 92.800 160.200 93.100 ;
        RECT 160.600 92.800 161.000 93.200 ;
        RECT 167.800 93.100 168.200 93.200 ;
        RECT 173.400 93.100 173.800 93.200 ;
        RECT 167.800 92.800 173.800 93.100 ;
        RECT 140.600 92.200 140.900 92.800 ;
        RECT 20.600 92.100 21.000 92.200 ;
        RECT 31.000 92.100 31.400 92.200 ;
        RECT 42.200 92.100 42.600 92.200 ;
        RECT 20.600 91.800 42.600 92.100 ;
        RECT 44.600 92.100 45.000 92.200 ;
        RECT 59.800 92.100 60.200 92.200 ;
        RECT 44.600 91.800 60.200 92.100 ;
        RECT 64.600 92.100 65.000 92.200 ;
        RECT 68.600 92.100 69.000 92.200 ;
        RECT 64.600 91.800 69.000 92.100 ;
        RECT 73.400 92.100 73.800 92.200 ;
        RECT 80.600 92.100 81.000 92.200 ;
        RECT 115.800 92.100 116.200 92.200 ;
        RECT 73.400 91.800 116.200 92.100 ;
        RECT 125.400 92.100 125.800 92.200 ;
        RECT 134.200 92.100 134.600 92.200 ;
        RECT 125.400 91.800 134.600 92.100 ;
        RECT 140.600 91.800 141.000 92.200 ;
        RECT 161.400 92.100 161.800 92.200 ;
        RECT 141.400 91.800 161.800 92.100 ;
        RECT 171.800 92.100 172.200 92.200 ;
        RECT 178.200 92.100 178.600 92.200 ;
        RECT 192.600 92.100 193.000 92.200 ;
        RECT 171.800 91.800 193.000 92.100 ;
        RECT 21.400 91.100 21.800 91.200 ;
        RECT 27.800 91.100 28.200 91.200 ;
        RECT 21.400 90.800 28.200 91.100 ;
        RECT 29.400 91.100 29.800 91.200 ;
        RECT 37.400 91.100 37.800 91.200 ;
        RECT 55.800 91.100 56.200 91.200 ;
        RECT 29.400 90.800 56.200 91.100 ;
        RECT 61.400 91.100 61.800 91.200 ;
        RECT 67.000 91.100 67.400 91.200 ;
        RECT 61.400 90.800 67.400 91.100 ;
        RECT 72.600 91.100 73.000 91.200 ;
        RECT 75.800 91.100 76.200 91.200 ;
        RECT 72.600 90.800 76.200 91.100 ;
        RECT 85.400 91.100 85.800 91.200 ;
        RECT 88.600 91.100 89.000 91.200 ;
        RECT 85.400 90.800 89.000 91.100 ;
        RECT 104.600 91.100 105.000 91.200 ;
        RECT 137.400 91.100 137.800 91.200 ;
        RECT 141.400 91.100 141.700 91.800 ;
        RECT 104.600 90.800 141.700 91.100 ;
        RECT 150.200 91.100 150.600 91.200 ;
        RECT 159.800 91.100 160.200 91.200 ;
        RECT 177.400 91.100 177.800 91.200 ;
        RECT 150.200 90.800 177.800 91.100 ;
        RECT 15.000 90.100 15.400 90.200 ;
        RECT 19.800 90.100 20.200 90.200 ;
        RECT 15.000 89.800 20.200 90.100 ;
        RECT 30.200 90.100 30.600 90.200 ;
        RECT 31.000 90.100 31.400 90.200 ;
        RECT 34.200 90.100 34.600 90.200 ;
        RECT 37.400 90.100 37.800 90.200 ;
        RECT 43.000 90.100 43.400 90.200 ;
        RECT 66.200 90.100 66.600 90.200 ;
        RECT 30.200 89.800 66.600 90.100 ;
        RECT 82.200 90.100 82.600 90.200 ;
        RECT 87.000 90.100 87.400 90.200 ;
        RECT 125.400 90.100 125.800 90.200 ;
        RECT 82.200 89.800 87.400 90.100 ;
        RECT 103.800 89.800 125.800 90.100 ;
        RECT 130.200 90.100 130.600 90.200 ;
        RECT 131.800 90.100 132.200 90.200 ;
        RECT 133.400 90.100 133.800 90.200 ;
        RECT 130.200 89.800 133.800 90.100 ;
        RECT 147.000 90.100 147.400 90.200 ;
        RECT 158.200 90.100 158.600 90.200 ;
        RECT 147.000 89.800 158.600 90.100 ;
        RECT 163.800 90.100 164.200 90.200 ;
        RECT 174.200 90.100 174.600 90.200 ;
        RECT 178.200 90.100 178.600 90.200 ;
        RECT 163.800 89.800 178.600 90.100 ;
        RECT 15.000 89.100 15.400 89.200 ;
        RECT 17.400 89.100 17.800 89.200 ;
        RECT 15.000 88.800 17.800 89.100 ;
        RECT 25.400 89.100 25.800 89.200 ;
        RECT 32.600 89.100 33.000 89.200 ;
        RECT 25.400 88.800 33.000 89.100 ;
        RECT 37.400 88.800 37.800 89.200 ;
        RECT 43.800 89.100 44.200 89.200 ;
        RECT 45.400 89.100 45.800 89.200 ;
        RECT 43.800 88.800 45.800 89.100 ;
        RECT 50.200 89.100 50.600 89.200 ;
        RECT 59.000 89.100 59.400 89.200 ;
        RECT 50.200 88.800 59.400 89.100 ;
        RECT 60.600 89.100 61.000 89.200 ;
        RECT 63.800 89.100 64.200 89.200 ;
        RECT 65.400 89.100 65.800 89.200 ;
        RECT 70.200 89.100 70.600 89.200 ;
        RECT 60.600 88.800 70.600 89.100 ;
        RECT 71.800 89.100 72.200 89.200 ;
        RECT 74.200 89.100 74.600 89.200 ;
        RECT 71.800 88.800 74.600 89.100 ;
        RECT 83.000 89.100 83.400 89.200 ;
        RECT 83.800 89.100 84.200 89.200 ;
        RECT 83.000 88.800 84.200 89.100 ;
        RECT 84.600 89.100 85.000 89.200 ;
        RECT 85.400 89.100 85.800 89.200 ;
        RECT 84.600 88.800 85.800 89.100 ;
        RECT 90.200 89.100 90.600 89.200 ;
        RECT 103.800 89.100 104.100 89.800 ;
        RECT 90.200 88.800 104.100 89.100 ;
        RECT 104.600 89.100 105.000 89.200 ;
        RECT 105.400 89.100 105.800 89.200 ;
        RECT 104.600 88.800 105.800 89.100 ;
        RECT 115.000 89.100 115.400 89.200 ;
        RECT 115.800 89.100 116.200 89.200 ;
        RECT 115.000 88.800 116.200 89.100 ;
        RECT 135.000 89.100 135.400 89.200 ;
        RECT 147.800 89.100 148.200 89.200 ;
        RECT 150.200 89.100 150.600 89.200 ;
        RECT 135.000 88.800 150.600 89.100 ;
        RECT 151.800 89.100 152.200 89.200 ;
        RECT 159.000 89.100 159.400 89.200 ;
        RECT 151.800 88.800 159.400 89.100 ;
        RECT 159.800 89.100 160.200 89.200 ;
        RECT 164.600 89.100 165.000 89.200 ;
        RECT 159.800 88.800 165.000 89.100 ;
        RECT 175.800 89.100 176.200 89.200 ;
        RECT 176.600 89.100 177.000 89.200 ;
        RECT 179.000 89.100 179.400 89.200 ;
        RECT 175.800 88.800 179.400 89.100 ;
        RECT 0.600 88.100 1.000 88.200 ;
        RECT 10.200 88.100 10.600 88.200 ;
        RECT 18.200 88.100 18.600 88.200 ;
        RECT 0.600 87.800 18.600 88.100 ;
        RECT 19.000 88.100 19.400 88.200 ;
        RECT 23.000 88.100 23.400 88.200 ;
        RECT 19.000 87.800 23.400 88.100 ;
        RECT 25.400 87.800 25.800 88.200 ;
        RECT 27.800 88.100 28.200 88.200 ;
        RECT 37.400 88.100 37.700 88.800 ;
        RECT 27.800 87.800 37.700 88.100 ;
        RECT 43.800 88.100 44.200 88.200 ;
        RECT 63.000 88.100 63.400 88.200 ;
        RECT 65.400 88.100 65.800 88.200 ;
        RECT 100.600 88.100 101.000 88.200 ;
        RECT 43.800 87.800 62.500 88.100 ;
        RECT 63.000 87.800 101.000 88.100 ;
        RECT 103.800 88.100 104.200 88.200 ;
        RECT 136.600 88.100 137.000 88.200 ;
        RECT 103.800 87.800 137.000 88.100 ;
        RECT 142.200 88.100 142.600 88.200 ;
        RECT 165.400 88.100 165.800 88.200 ;
        RECT 142.200 87.800 165.800 88.100 ;
        RECT 179.000 88.100 179.400 88.200 ;
        RECT 196.600 88.100 197.000 88.200 ;
        RECT 179.000 87.800 197.000 88.100 ;
        RECT 7.000 86.800 7.400 87.200 ;
        RECT 8.600 87.100 9.000 87.200 ;
        RECT 25.400 87.100 25.700 87.800 ;
        RECT 8.600 86.800 25.700 87.100 ;
        RECT 35.800 87.100 36.200 87.200 ;
        RECT 39.000 87.100 39.400 87.200 ;
        RECT 44.600 87.100 45.000 87.200 ;
        RECT 35.800 86.800 45.000 87.100 ;
        RECT 62.200 87.100 62.500 87.800 ;
        RECT 75.000 87.100 75.400 87.200 ;
        RECT 62.200 86.800 75.400 87.100 ;
        RECT 79.800 86.800 80.200 87.200 ;
        RECT 83.000 87.100 83.400 87.200 ;
        RECT 87.800 87.100 88.200 87.200 ;
        RECT 83.000 86.800 88.200 87.100 ;
        RECT 92.600 87.100 93.000 87.200 ;
        RECT 99.000 87.100 99.400 87.200 ;
        RECT 92.600 86.800 99.400 87.100 ;
        RECT 106.200 86.800 106.600 87.200 ;
        RECT 122.200 87.100 122.600 87.200 ;
        RECT 114.200 86.800 122.600 87.100 ;
        RECT 125.400 87.100 125.800 87.200 ;
        RECT 131.800 87.100 132.200 87.200 ;
        RECT 125.400 86.800 132.200 87.100 ;
        RECT 143.800 86.800 144.200 87.200 ;
        RECT 164.600 87.100 165.000 87.200 ;
        RECT 145.400 86.800 165.000 87.100 ;
        RECT 170.200 87.100 170.600 87.200 ;
        RECT 176.600 87.100 177.000 87.200 ;
        RECT 179.000 87.100 179.300 87.800 ;
        RECT 170.200 86.800 171.300 87.100 ;
        RECT 176.600 86.800 179.300 87.100 ;
        RECT 191.000 86.800 191.400 87.200 ;
        RECT 192.600 86.800 193.000 87.200 ;
        RECT 7.000 86.100 7.300 86.800 ;
        RECT 11.800 86.100 12.200 86.200 ;
        RECT 7.000 85.800 12.200 86.100 ;
        RECT 12.600 86.100 13.000 86.200 ;
        RECT 13.400 86.100 13.800 86.200 ;
        RECT 15.800 86.100 16.200 86.200 ;
        RECT 12.600 85.800 16.200 86.100 ;
        RECT 17.400 86.100 17.800 86.200 ;
        RECT 22.200 86.100 22.600 86.200 ;
        RECT 17.400 85.800 22.600 86.100 ;
        RECT 34.200 86.100 34.600 86.200 ;
        RECT 40.600 86.100 41.000 86.200 ;
        RECT 45.400 86.100 45.800 86.200 ;
        RECT 34.200 85.800 40.100 86.100 ;
        RECT 40.600 85.800 45.800 86.100 ;
        RECT 55.000 86.100 55.400 86.300 ;
        RECT 60.600 86.100 61.000 86.200 ;
        RECT 55.000 85.800 61.000 86.100 ;
        RECT 74.200 86.100 74.600 86.200 ;
        RECT 75.000 86.100 75.400 86.200 ;
        RECT 74.200 85.800 75.400 86.100 ;
        RECT 77.400 86.100 77.800 86.200 ;
        RECT 78.200 86.100 78.600 86.200 ;
        RECT 77.400 85.800 78.600 86.100 ;
        RECT 79.800 86.100 80.100 86.800 ;
        RECT 99.000 86.200 99.300 86.800 ;
        RECT 106.200 86.200 106.500 86.800 ;
        RECT 114.200 86.200 114.500 86.800 ;
        RECT 143.800 86.200 144.100 86.800 ;
        RECT 145.400 86.200 145.700 86.800 ;
        RECT 171.000 86.200 171.300 86.800 ;
        RECT 191.000 86.200 191.300 86.800 ;
        RECT 82.200 86.100 82.600 86.200 ;
        RECT 79.800 85.800 82.600 86.100 ;
        RECT 83.800 86.100 84.200 86.200 ;
        RECT 87.000 86.100 87.400 86.200 ;
        RECT 83.800 85.800 87.400 86.100 ;
        RECT 99.000 85.800 99.400 86.200 ;
        RECT 100.600 86.100 101.000 86.200 ;
        RECT 103.800 86.100 104.200 86.200 ;
        RECT 100.600 85.800 104.200 86.100 ;
        RECT 106.200 85.800 106.600 86.200 ;
        RECT 114.200 85.800 114.600 86.200 ;
        RECT 119.000 86.100 119.400 86.200 ;
        RECT 128.600 86.100 129.000 86.200 ;
        RECT 119.000 85.800 129.000 86.100 ;
        RECT 143.800 85.800 144.200 86.200 ;
        RECT 145.400 85.800 145.800 86.200 ;
        RECT 149.400 86.100 149.800 86.200 ;
        RECT 151.800 86.100 152.200 86.200 ;
        RECT 149.400 85.800 152.200 86.100 ;
        RECT 156.600 86.100 157.000 86.200 ;
        RECT 166.200 86.100 166.600 86.200 ;
        RECT 156.600 85.800 166.600 86.100 ;
        RECT 171.000 85.800 171.400 86.200 ;
        RECT 177.400 86.100 177.800 86.200 ;
        RECT 184.600 86.100 185.000 86.200 ;
        RECT 177.400 85.800 185.000 86.100 ;
        RECT 191.000 85.800 191.400 86.200 ;
        RECT 192.600 86.100 192.900 86.800 ;
        RECT 195.000 86.100 195.400 86.200 ;
        RECT 192.600 85.800 195.400 86.100 ;
        RECT 200.600 86.100 201.000 86.200 ;
        RECT 201.400 86.100 201.800 86.200 ;
        RECT 200.600 85.800 201.800 86.100 ;
        RECT 39.800 85.200 40.100 85.800 ;
        RECT 100.600 85.200 100.900 85.800 ;
        RECT 39.800 84.800 40.200 85.200 ;
        RECT 61.400 85.100 61.800 85.200 ;
        RECT 63.000 85.100 63.400 85.200 ;
        RECT 61.400 84.800 63.400 85.100 ;
        RECT 68.600 85.100 69.000 85.200 ;
        RECT 71.800 85.100 72.200 85.200 ;
        RECT 79.000 85.100 79.400 85.200 ;
        RECT 80.600 85.100 81.000 85.200 ;
        RECT 68.600 84.800 78.500 85.100 ;
        RECT 79.000 84.800 81.000 85.100 ;
        RECT 100.600 84.800 101.000 85.200 ;
        RECT 103.000 85.100 103.400 85.200 ;
        RECT 110.200 85.100 110.600 85.200 ;
        RECT 103.000 84.800 110.600 85.100 ;
        RECT 116.600 85.100 117.000 85.200 ;
        RECT 147.800 85.100 148.200 85.200 ;
        RECT 116.600 84.800 148.200 85.100 ;
        RECT 159.000 85.100 159.400 85.200 ;
        RECT 162.200 85.100 162.600 85.200 ;
        RECT 159.000 84.800 162.600 85.100 ;
        RECT 166.200 85.100 166.600 85.200 ;
        RECT 171.000 85.100 171.400 85.200 ;
        RECT 185.400 85.100 185.800 85.200 ;
        RECT 191.800 85.100 192.200 85.200 ;
        RECT 193.400 85.100 193.800 85.200 ;
        RECT 166.200 84.800 172.100 85.100 ;
        RECT 185.400 84.800 193.800 85.100 ;
        RECT 78.200 84.200 78.500 84.800 ;
        RECT 39.000 84.100 39.400 84.200 ;
        RECT 60.600 84.100 61.000 84.200 ;
        RECT 39.000 83.800 61.000 84.100 ;
        RECT 72.600 83.800 73.000 84.200 ;
        RECT 78.200 83.800 78.600 84.200 ;
        RECT 86.200 84.100 86.600 84.200 ;
        RECT 91.000 84.100 91.400 84.200 ;
        RECT 96.600 84.100 97.000 84.200 ;
        RECT 147.000 84.100 147.400 84.200 ;
        RECT 159.000 84.100 159.400 84.200 ;
        RECT 171.000 84.100 171.400 84.200 ;
        RECT 86.200 83.800 171.400 84.100 ;
        RECT 172.600 84.100 173.000 84.200 ;
        RECT 191.000 84.100 191.400 84.200 ;
        RECT 172.600 83.800 191.400 84.100 ;
        RECT 15.800 83.100 16.200 83.200 ;
        RECT 18.200 83.100 18.600 83.200 ;
        RECT 58.200 83.100 58.600 83.200 ;
        RECT 15.800 82.800 58.600 83.100 ;
        RECT 62.200 83.100 62.600 83.200 ;
        RECT 64.600 83.100 65.000 83.200 ;
        RECT 62.200 82.800 65.000 83.100 ;
        RECT 65.400 83.100 65.800 83.200 ;
        RECT 72.600 83.100 72.900 83.800 ;
        RECT 65.400 82.800 72.900 83.100 ;
        RECT 83.000 83.100 83.400 83.200 ;
        RECT 115.800 83.100 116.200 83.200 ;
        RECT 83.000 82.800 116.200 83.100 ;
        RECT 133.400 83.100 133.800 83.200 ;
        RECT 153.400 83.100 153.800 83.200 ;
        RECT 168.600 83.100 169.000 83.200 ;
        RECT 190.200 83.100 190.600 83.200 ;
        RECT 203.800 83.100 204.200 83.200 ;
        RECT 133.400 82.800 204.200 83.100 ;
        RECT 9.400 82.100 9.800 82.200 ;
        RECT 41.400 82.100 41.800 82.200 ;
        RECT 9.400 81.800 41.800 82.100 ;
        RECT 52.600 82.100 53.000 82.200 ;
        RECT 58.200 82.100 58.600 82.200 ;
        RECT 52.600 81.800 58.600 82.100 ;
        RECT 61.400 82.100 61.800 82.200 ;
        RECT 91.800 82.100 92.200 82.200 ;
        RECT 61.400 81.800 92.200 82.100 ;
        RECT 94.200 82.100 94.600 82.200 ;
        RECT 95.000 82.100 95.400 82.200 ;
        RECT 94.200 81.800 95.400 82.100 ;
        RECT 163.000 81.800 163.400 82.200 ;
        RECT 163.000 81.200 163.300 81.800 ;
        RECT 11.800 81.100 12.200 81.200 ;
        RECT 13.400 81.100 13.800 81.200 ;
        RECT 14.200 81.100 14.600 81.200 ;
        RECT 18.200 81.100 18.600 81.200 ;
        RECT 47.000 81.100 47.400 81.200 ;
        RECT 11.800 80.800 47.400 81.100 ;
        RECT 70.200 81.100 70.600 81.200 ;
        RECT 72.600 81.100 73.000 81.200 ;
        RECT 70.200 80.800 73.000 81.100 ;
        RECT 83.000 81.100 83.400 81.200 ;
        RECT 94.200 81.100 94.600 81.200 ;
        RECT 83.000 80.800 94.600 81.100 ;
        RECT 163.000 80.800 163.400 81.200 ;
        RECT 23.800 80.100 24.200 80.200 ;
        RECT 31.000 80.100 31.400 80.200 ;
        RECT 23.800 79.800 31.400 80.100 ;
        RECT 42.200 80.100 42.600 80.200 ;
        RECT 47.800 80.100 48.200 80.200 ;
        RECT 42.200 79.800 48.200 80.100 ;
        RECT 95.800 80.100 96.200 80.200 ;
        RECT 97.400 80.100 97.800 80.200 ;
        RECT 95.800 79.800 97.800 80.100 ;
        RECT 22.200 79.100 22.600 79.200 ;
        RECT 27.000 79.100 27.400 79.200 ;
        RECT 22.200 78.800 27.400 79.100 ;
        RECT 45.400 79.100 45.800 79.200 ;
        RECT 50.200 79.100 50.600 79.200 ;
        RECT 45.400 78.800 50.600 79.100 ;
        RECT 53.400 78.800 53.800 79.200 ;
        RECT 76.600 79.100 77.000 79.200 ;
        RECT 77.400 79.100 77.800 79.200 ;
        RECT 76.600 78.800 77.800 79.100 ;
        RECT 80.600 79.100 81.000 79.200 ;
        RECT 115.000 79.100 115.400 79.200 ;
        RECT 80.600 78.800 115.400 79.100 ;
        RECT 115.800 79.100 116.200 79.200 ;
        RECT 119.000 79.100 119.400 79.200 ;
        RECT 115.800 78.800 119.400 79.100 ;
        RECT 148.600 79.100 149.000 79.200 ;
        RECT 153.400 79.100 153.800 79.200 ;
        RECT 148.600 78.800 153.800 79.100 ;
        RECT 42.200 78.100 42.600 78.200 ;
        RECT 52.600 78.100 53.000 78.200 ;
        RECT 42.200 77.800 53.000 78.100 ;
        RECT 53.400 78.100 53.700 78.800 ;
        RECT 61.400 78.100 61.800 78.200 ;
        RECT 53.400 77.800 61.800 78.100 ;
        RECT 69.400 78.100 69.800 78.200 ;
        RECT 86.200 78.100 86.600 78.200 ;
        RECT 99.800 78.100 100.200 78.200 ;
        RECT 100.600 78.100 101.000 78.200 ;
        RECT 118.200 78.100 118.600 78.200 ;
        RECT 69.400 77.800 118.600 78.100 ;
        RECT 119.000 78.100 119.400 78.200 ;
        RECT 167.800 78.100 168.200 78.200 ;
        RECT 119.000 77.800 168.200 78.100 ;
        RECT 30.200 77.100 30.600 77.200 ;
        RECT 39.800 77.100 40.200 77.200 ;
        RECT 52.600 77.100 53.000 77.200 ;
        RECT 30.200 76.800 53.000 77.100 ;
        RECT 55.000 76.800 55.400 77.200 ;
        RECT 72.600 77.100 73.000 77.200 ;
        RECT 83.800 77.100 84.200 77.200 ;
        RECT 72.600 76.800 84.200 77.100 ;
        RECT 91.800 77.100 92.200 77.200 ;
        RECT 93.400 77.100 93.800 77.200 ;
        RECT 91.800 76.800 93.800 77.100 ;
        RECT 95.800 77.100 96.200 77.200 ;
        RECT 99.000 77.100 99.400 77.200 ;
        RECT 95.800 76.800 99.400 77.100 ;
        RECT 119.800 77.100 120.200 77.200 ;
        RECT 131.000 77.100 131.400 77.200 ;
        RECT 119.800 76.800 131.400 77.100 ;
        RECT 137.400 77.100 137.800 77.200 ;
        RECT 139.800 77.100 140.200 77.200 ;
        RECT 140.600 77.100 141.000 77.200 ;
        RECT 137.400 76.800 141.000 77.100 ;
        RECT 141.400 77.100 141.800 77.200 ;
        RECT 150.200 77.100 150.600 77.200 ;
        RECT 156.600 77.100 157.000 77.200 ;
        RECT 141.400 76.800 157.000 77.100 ;
        RECT 160.600 77.100 161.000 77.200 ;
        RECT 172.600 77.100 173.000 77.200 ;
        RECT 160.600 76.800 173.000 77.100 ;
        RECT 175.800 77.100 176.200 77.200 ;
        RECT 175.800 76.800 181.700 77.100 ;
        RECT 21.400 75.800 21.800 76.200 ;
        RECT 44.600 76.100 45.000 76.200 ;
        RECT 47.000 76.100 47.400 76.200 ;
        RECT 44.600 75.800 47.400 76.100 ;
        RECT 48.600 76.100 49.000 76.200 ;
        RECT 49.400 76.100 49.800 76.200 ;
        RECT 48.600 75.800 49.800 76.100 ;
        RECT 51.000 76.100 51.400 76.200 ;
        RECT 54.200 76.100 54.600 76.200 ;
        RECT 55.000 76.100 55.300 76.800 ;
        RECT 181.400 76.200 181.700 76.800 ;
        RECT 51.000 75.800 55.300 76.100 ;
        RECT 67.800 76.100 68.200 76.200 ;
        RECT 70.200 76.100 70.600 76.200 ;
        RECT 67.800 75.800 70.600 76.100 ;
        RECT 71.000 76.100 71.400 76.200 ;
        RECT 71.800 76.100 72.200 76.200 ;
        RECT 71.000 75.800 72.200 76.100 ;
        RECT 75.000 76.100 75.400 76.200 ;
        RECT 87.800 76.100 88.200 76.200 ;
        RECT 75.000 75.800 88.200 76.100 ;
        RECT 88.600 76.100 89.000 76.200 ;
        RECT 97.400 76.100 97.800 76.200 ;
        RECT 88.600 75.800 97.800 76.100 ;
        RECT 104.600 76.100 105.000 76.200 ;
        RECT 107.000 76.100 107.400 76.200 ;
        RECT 108.600 76.100 109.000 76.200 ;
        RECT 111.800 76.100 112.200 76.200 ;
        RECT 104.600 75.800 112.200 76.100 ;
        RECT 113.400 76.100 113.800 76.200 ;
        RECT 115.000 76.100 115.400 76.200 ;
        RECT 113.400 75.800 115.400 76.100 ;
        RECT 132.600 76.100 133.000 76.200 ;
        RECT 135.000 76.100 135.400 76.200 ;
        RECT 132.600 75.800 135.400 76.100 ;
        RECT 135.800 76.100 136.200 76.200 ;
        RECT 147.800 76.100 148.200 76.200 ;
        RECT 135.800 75.800 148.200 76.100 ;
        RECT 149.400 76.100 149.800 76.200 ;
        RECT 157.400 76.100 157.800 76.200 ;
        RECT 149.400 75.800 157.800 76.100 ;
        RECT 158.200 76.100 158.600 76.200 ;
        RECT 159.000 76.100 159.400 76.200 ;
        RECT 158.200 75.800 159.400 76.100 ;
        RECT 160.600 76.100 161.000 76.200 ;
        RECT 161.400 76.100 161.800 76.200 ;
        RECT 160.600 75.800 161.800 76.100 ;
        RECT 165.400 76.100 165.800 76.200 ;
        RECT 167.800 76.100 168.200 76.200 ;
        RECT 165.400 75.800 168.200 76.100 ;
        RECT 181.400 75.800 181.800 76.200 ;
        RECT 5.400 75.100 5.800 75.200 ;
        RECT 13.400 75.100 13.800 75.200 ;
        RECT 5.400 74.800 13.800 75.100 ;
        RECT 14.200 74.800 14.600 75.200 ;
        RECT 16.600 75.100 17.000 75.200 ;
        RECT 21.400 75.100 21.700 75.800 ;
        RECT 47.000 75.200 47.300 75.800 ;
        RECT 16.600 74.800 21.700 75.100 ;
        RECT 33.400 74.800 33.800 75.200 ;
        RECT 36.600 75.100 37.000 75.200 ;
        RECT 43.800 75.100 44.200 75.200 ;
        RECT 36.600 74.800 44.200 75.100 ;
        RECT 47.000 74.800 47.400 75.200 ;
        RECT 47.800 75.100 48.200 75.200 ;
        RECT 51.000 75.100 51.400 75.200 ;
        RECT 55.000 75.100 55.400 75.200 ;
        RECT 47.800 74.800 55.400 75.100 ;
        RECT 59.000 74.800 59.400 75.200 ;
        RECT 60.600 75.100 61.000 75.200 ;
        RECT 60.600 74.800 62.500 75.100 ;
        RECT 14.200 74.200 14.500 74.800 ;
        RECT 11.800 74.100 12.200 74.200 ;
        RECT 14.200 74.100 14.600 74.200 ;
        RECT 18.200 74.100 18.600 74.200 ;
        RECT 11.800 73.800 18.600 74.100 ;
        RECT 24.600 74.100 25.000 74.200 ;
        RECT 33.400 74.100 33.700 74.800 ;
        RECT 59.000 74.200 59.300 74.800 ;
        RECT 62.200 74.200 62.500 74.800 ;
        RECT 63.000 74.800 63.400 75.200 ;
        RECT 66.200 75.100 66.600 75.200 ;
        RECT 67.000 75.100 67.400 75.200 ;
        RECT 66.200 74.800 67.400 75.100 ;
        RECT 72.600 75.100 73.000 75.200 ;
        RECT 73.400 75.100 73.800 75.200 ;
        RECT 72.600 74.800 73.800 75.100 ;
        RECT 74.200 75.100 74.600 75.200 ;
        RECT 75.000 75.100 75.400 75.200 ;
        RECT 74.200 74.800 75.400 75.100 ;
        RECT 75.800 75.100 76.200 75.200 ;
        RECT 76.600 75.100 77.000 75.200 ;
        RECT 75.800 74.800 77.000 75.100 ;
        RECT 79.000 75.100 79.400 75.200 ;
        RECT 84.600 75.100 85.000 75.200 ;
        RECT 79.000 74.800 85.000 75.100 ;
        RECT 88.600 75.100 89.000 75.200 ;
        RECT 93.400 75.100 93.800 75.200 ;
        RECT 88.600 74.800 93.800 75.100 ;
        RECT 96.600 75.100 97.000 75.200 ;
        RECT 105.400 75.100 105.800 75.200 ;
        RECT 96.600 74.800 105.800 75.100 ;
        RECT 106.200 75.100 106.600 75.200 ;
        RECT 116.600 75.100 117.000 75.200 ;
        RECT 129.400 75.100 129.800 75.200 ;
        RECT 106.200 74.800 117.000 75.100 ;
        RECT 124.600 74.800 129.800 75.100 ;
        RECT 130.200 75.100 130.600 75.200 ;
        RECT 159.800 75.100 160.200 75.200 ;
        RECT 176.600 75.100 177.000 75.200 ;
        RECT 179.800 75.100 180.200 75.200 ;
        RECT 130.200 74.800 180.200 75.100 ;
        RECT 194.200 74.800 194.600 75.200 ;
        RECT 195.800 75.100 196.200 75.200 ;
        RECT 199.800 75.100 200.200 75.200 ;
        RECT 195.800 74.800 200.200 75.100 ;
        RECT 24.600 73.800 33.700 74.100 ;
        RECT 46.200 74.100 46.600 74.200 ;
        RECT 53.400 74.100 53.800 74.200 ;
        RECT 46.200 73.800 53.800 74.100 ;
        RECT 59.000 73.800 59.400 74.200 ;
        RECT 62.200 73.800 62.600 74.200 ;
        RECT 63.000 74.100 63.300 74.800 ;
        RECT 124.600 74.700 125.000 74.800 ;
        RECT 194.200 74.200 194.500 74.800 ;
        RECT 66.200 74.100 66.600 74.200 ;
        RECT 63.000 73.800 66.600 74.100 ;
        RECT 67.000 74.100 67.400 74.200 ;
        RECT 67.800 74.100 68.200 74.200 ;
        RECT 67.000 73.800 68.200 74.100 ;
        RECT 71.000 74.100 71.400 74.200 ;
        RECT 73.400 74.100 73.800 74.200 ;
        RECT 71.000 73.800 73.800 74.100 ;
        RECT 75.000 74.100 75.400 74.200 ;
        RECT 77.400 74.100 77.800 74.200 ;
        RECT 78.200 74.100 78.600 74.200 ;
        RECT 75.000 73.800 76.100 74.100 ;
        RECT 77.400 73.800 78.600 74.100 ;
        RECT 82.200 74.100 82.600 74.200 ;
        RECT 83.000 74.100 83.400 74.200 ;
        RECT 82.200 73.800 83.400 74.100 ;
        RECT 83.800 74.100 84.200 74.200 ;
        RECT 89.400 74.100 89.800 74.200 ;
        RECT 83.800 73.800 89.800 74.100 ;
        RECT 91.000 74.100 91.400 74.200 ;
        RECT 91.800 74.100 92.200 74.200 ;
        RECT 91.000 73.800 92.200 74.100 ;
        RECT 97.400 74.100 97.800 74.200 ;
        RECT 107.000 74.100 107.400 74.200 ;
        RECT 97.400 73.800 107.400 74.100 ;
        RECT 112.600 74.100 113.000 74.200 ;
        RECT 123.800 74.100 124.200 74.200 ;
        RECT 112.600 73.800 124.200 74.100 ;
        RECT 124.600 74.100 125.000 74.200 ;
        RECT 143.800 74.100 144.200 74.200 ;
        RECT 144.600 74.100 145.000 74.200 ;
        RECT 124.600 73.800 143.300 74.100 ;
        RECT 143.800 73.800 145.000 74.100 ;
        RECT 154.200 74.100 154.600 74.200 ;
        RECT 155.000 74.100 155.400 74.200 ;
        RECT 158.200 74.100 158.600 74.200 ;
        RECT 159.800 74.100 160.200 74.200 ;
        RECT 154.200 73.800 155.400 74.100 ;
        RECT 157.400 73.800 160.200 74.100 ;
        RECT 160.600 74.100 161.000 74.200 ;
        RECT 170.200 74.100 170.600 74.200 ;
        RECT 173.400 74.100 173.800 74.200 ;
        RECT 160.600 73.800 173.800 74.100 ;
        RECT 179.000 74.100 179.400 74.200 ;
        RECT 186.200 74.100 186.600 74.200 ;
        RECT 179.000 73.800 186.600 74.100 ;
        RECT 191.800 73.800 192.200 74.200 ;
        RECT 194.200 74.100 194.600 74.200 ;
        RECT 199.800 74.100 200.200 74.200 ;
        RECT 194.200 73.800 200.200 74.100 ;
        RECT 75.800 73.200 76.100 73.800 ;
        RECT 143.000 73.200 143.300 73.800 ;
        RECT 17.400 73.100 17.800 73.200 ;
        RECT 18.200 73.100 18.600 73.200 ;
        RECT 35.000 73.100 35.400 73.200 ;
        RECT 17.400 72.800 18.600 73.100 ;
        RECT 31.800 72.800 35.400 73.100 ;
        RECT 43.800 73.100 44.200 73.200 ;
        RECT 47.800 73.100 48.200 73.200 ;
        RECT 68.600 73.100 69.000 73.200 ;
        RECT 71.800 73.100 72.200 73.200 ;
        RECT 43.800 72.800 48.200 73.100 ;
        RECT 67.800 72.800 72.200 73.100 ;
        RECT 75.800 72.800 76.200 73.200 ;
        RECT 78.200 73.100 78.600 73.200 ;
        RECT 79.800 73.100 80.200 73.200 ;
        RECT 78.200 72.800 80.200 73.100 ;
        RECT 80.600 73.100 81.000 73.200 ;
        RECT 83.000 73.100 83.400 73.200 ;
        RECT 80.600 72.800 83.400 73.100 ;
        RECT 84.600 73.100 85.000 73.200 ;
        RECT 95.000 73.100 95.400 73.200 ;
        RECT 84.600 72.800 95.400 73.100 ;
        RECT 102.200 73.100 102.600 73.200 ;
        RECT 109.400 73.100 109.800 73.200 ;
        RECT 102.200 72.800 109.800 73.100 ;
        RECT 111.000 73.100 111.400 73.200 ;
        RECT 113.400 73.100 113.800 73.200 ;
        RECT 111.000 72.800 113.800 73.100 ;
        RECT 115.000 73.100 115.400 73.200 ;
        RECT 115.800 73.100 116.200 73.200 ;
        RECT 128.600 73.100 129.000 73.200 ;
        RECT 115.000 72.800 129.000 73.100 ;
        RECT 129.400 73.100 129.800 73.200 ;
        RECT 135.000 73.100 135.400 73.200 ;
        RECT 139.800 73.100 140.200 73.200 ;
        RECT 142.200 73.100 142.600 73.200 ;
        RECT 129.400 72.800 135.400 73.100 ;
        RECT 139.000 72.800 142.600 73.100 ;
        RECT 143.000 72.800 143.400 73.200 ;
        RECT 144.600 73.100 145.000 73.200 ;
        RECT 154.200 73.100 154.600 73.200 ;
        RECT 163.800 73.100 164.200 73.200 ;
        RECT 169.400 73.100 169.800 73.200 ;
        RECT 144.600 72.800 155.300 73.100 ;
        RECT 163.800 72.800 169.800 73.100 ;
        RECT 191.800 73.100 192.100 73.800 ;
        RECT 193.400 73.100 193.800 73.200 ;
        RECT 191.800 72.800 193.800 73.100 ;
        RECT 195.800 73.100 196.200 73.200 ;
        RECT 199.000 73.100 199.400 73.200 ;
        RECT 195.800 72.800 199.400 73.100 ;
        RECT 31.800 72.200 32.100 72.800 ;
        RECT 31.800 71.800 32.200 72.200 ;
        RECT 32.600 72.100 33.000 72.200 ;
        RECT 60.600 72.100 61.000 72.200 ;
        RECT 69.400 72.100 69.800 72.200 ;
        RECT 32.600 71.800 69.800 72.100 ;
        RECT 85.400 72.100 85.800 72.200 ;
        RECT 88.600 72.100 89.000 72.200 ;
        RECT 85.400 71.800 89.000 72.100 ;
        RECT 90.200 72.100 90.600 72.200 ;
        RECT 116.600 72.100 117.000 72.200 ;
        RECT 122.200 72.100 122.600 72.200 ;
        RECT 90.200 71.800 122.600 72.100 ;
        RECT 136.600 72.100 137.000 72.200 ;
        RECT 168.600 72.100 169.000 72.200 ;
        RECT 180.600 72.100 181.000 72.200 ;
        RECT 136.600 71.800 181.000 72.100 ;
        RECT 15.000 71.100 15.400 71.200 ;
        RECT 28.600 71.100 29.000 71.200 ;
        RECT 15.000 70.800 29.000 71.100 ;
        RECT 51.800 71.100 52.200 71.200 ;
        RECT 87.800 71.100 88.200 71.200 ;
        RECT 51.800 70.800 88.200 71.100 ;
        RECT 181.400 71.100 181.800 71.200 ;
        RECT 184.600 71.100 185.000 71.200 ;
        RECT 181.400 70.800 185.000 71.100 ;
        RECT 24.600 70.100 25.000 70.200 ;
        RECT 28.600 70.100 29.000 70.200 ;
        RECT 24.600 69.800 29.000 70.100 ;
        RECT 46.200 70.100 46.600 70.200 ;
        RECT 56.600 70.100 57.000 70.200 ;
        RECT 46.200 69.800 57.000 70.100 ;
        RECT 58.200 70.100 58.600 70.200 ;
        RECT 75.800 70.100 76.200 70.200 ;
        RECT 79.000 70.100 79.400 70.200 ;
        RECT 58.200 69.800 72.100 70.100 ;
        RECT 75.800 69.800 79.400 70.100 ;
        RECT 106.200 70.100 106.600 70.200 ;
        RECT 139.800 70.100 140.200 70.200 ;
        RECT 106.200 69.800 140.200 70.100 ;
        RECT 141.400 70.100 141.800 70.200 ;
        RECT 151.000 70.100 151.400 70.200 ;
        RECT 141.400 69.800 151.400 70.100 ;
        RECT 180.600 70.100 181.000 70.200 ;
        RECT 182.200 70.100 182.600 70.200 ;
        RECT 180.600 69.800 182.600 70.100 ;
        RECT 187.000 70.100 187.400 70.200 ;
        RECT 197.400 70.100 197.800 70.200 ;
        RECT 187.000 69.800 197.800 70.100 ;
        RECT 10.200 69.100 10.600 69.200 ;
        RECT 15.000 69.100 15.400 69.200 ;
        RECT 48.600 69.100 49.000 69.200 ;
        RECT 10.200 68.800 49.000 69.100 ;
        RECT 57.400 69.100 57.800 69.200 ;
        RECT 59.000 69.100 59.400 69.200 ;
        RECT 57.400 68.800 59.400 69.100 ;
        RECT 65.400 69.100 65.800 69.200 ;
        RECT 71.000 69.100 71.400 69.200 ;
        RECT 65.400 68.800 71.400 69.100 ;
        RECT 71.800 69.100 72.100 69.800 ;
        RECT 75.800 69.100 76.200 69.200 ;
        RECT 87.000 69.100 87.400 69.200 ;
        RECT 71.800 68.800 87.400 69.100 ;
        RECT 98.200 69.100 98.600 69.200 ;
        RECT 99.000 69.100 99.400 69.200 ;
        RECT 98.200 68.800 99.400 69.100 ;
        RECT 118.200 68.800 118.600 69.200 ;
        RECT 140.600 68.800 141.000 69.200 ;
        RECT 154.200 69.100 154.600 69.200 ;
        RECT 161.400 69.100 161.800 69.200 ;
        RECT 154.200 68.800 161.800 69.100 ;
        RECT 187.800 68.800 188.200 69.200 ;
        RECT 200.600 69.100 201.000 69.200 ;
        RECT 195.000 68.800 201.000 69.100 ;
        RECT 19.000 68.100 19.400 68.200 ;
        RECT 27.000 68.100 27.400 68.200 ;
        RECT 19.000 67.800 27.400 68.100 ;
        RECT 27.800 68.100 28.200 68.200 ;
        RECT 29.400 68.100 29.800 68.200 ;
        RECT 27.800 67.800 29.800 68.100 ;
        RECT 33.400 67.800 33.800 68.200 ;
        RECT 46.200 68.100 46.600 68.200 ;
        RECT 47.800 68.100 48.200 68.200 ;
        RECT 50.200 68.100 50.600 68.200 ;
        RECT 59.000 68.100 59.400 68.200 ;
        RECT 64.600 68.100 65.000 68.200 ;
        RECT 70.200 68.100 70.600 68.200 ;
        RECT 72.600 68.100 73.000 68.200 ;
        RECT 46.200 67.800 48.900 68.100 ;
        RECT 50.200 67.800 55.300 68.100 ;
        RECT 59.000 67.800 65.000 68.100 ;
        RECT 69.400 67.800 73.000 68.100 ;
        RECT 87.000 68.100 87.400 68.200 ;
        RECT 118.200 68.100 118.500 68.800 ;
        RECT 87.000 67.800 118.500 68.100 ;
        RECT 119.000 68.100 119.400 68.200 ;
        RECT 119.800 68.100 120.200 68.200 ;
        RECT 132.600 68.100 133.000 68.200 ;
        RECT 119.000 67.800 120.200 68.100 ;
        RECT 123.000 67.800 133.000 68.100 ;
        RECT 134.200 68.100 134.600 68.200 ;
        RECT 135.000 68.100 135.400 68.200 ;
        RECT 134.200 67.800 135.400 68.100 ;
        RECT 140.600 68.100 140.900 68.800 ;
        RECT 145.400 68.100 145.800 68.200 ;
        RECT 140.600 67.800 145.800 68.100 ;
        RECT 146.200 68.100 146.600 68.200 ;
        RECT 147.000 68.100 147.400 68.200 ;
        RECT 146.200 67.800 147.400 68.100 ;
        RECT 147.800 68.100 148.200 68.200 ;
        RECT 160.600 68.100 161.000 68.200 ;
        RECT 147.800 67.800 161.000 68.100 ;
        RECT 167.800 68.100 168.200 68.200 ;
        RECT 187.800 68.100 188.100 68.800 ;
        RECT 167.800 67.800 188.100 68.100 ;
        RECT 195.000 68.200 195.300 68.800 ;
        RECT 201.400 68.200 201.700 69.100 ;
        RECT 195.000 67.800 195.400 68.200 ;
        RECT 196.600 68.100 197.000 68.200 ;
        RECT 199.000 68.100 199.400 68.200 ;
        RECT 196.600 67.800 199.400 68.100 ;
        RECT 201.400 67.800 201.800 68.200 ;
        RECT 10.200 67.100 10.600 67.200 ;
        RECT 14.200 67.100 14.600 67.200 ;
        RECT 10.200 66.800 14.600 67.100 ;
        RECT 26.200 67.100 26.600 67.200 ;
        RECT 30.200 67.100 30.600 67.200 ;
        RECT 26.200 66.800 30.600 67.100 ;
        RECT 33.400 67.100 33.700 67.800 ;
        RECT 55.000 67.200 55.300 67.800 ;
        RECT 123.000 67.200 123.300 67.800 ;
        RECT 42.200 67.100 42.600 67.200 ;
        RECT 47.000 67.100 47.400 67.200 ;
        RECT 33.400 66.800 47.400 67.100 ;
        RECT 48.600 67.100 49.000 67.200 ;
        RECT 51.000 67.100 51.400 67.200 ;
        RECT 48.600 66.800 51.400 67.100 ;
        RECT 51.800 67.100 52.200 67.200 ;
        RECT 52.600 67.100 53.000 67.200 ;
        RECT 51.800 66.800 53.000 67.100 ;
        RECT 55.000 66.800 55.400 67.200 ;
        RECT 63.800 67.100 64.200 67.200 ;
        RECT 70.200 67.100 70.600 67.200 ;
        RECT 75.000 67.100 75.400 67.200 ;
        RECT 63.800 66.800 75.400 67.100 ;
        RECT 84.600 67.100 85.000 67.200 ;
        RECT 85.400 67.100 85.800 67.200 ;
        RECT 84.600 66.800 85.800 67.100 ;
        RECT 92.600 67.100 93.000 67.200 ;
        RECT 93.400 67.100 93.800 67.200 ;
        RECT 92.600 66.800 93.800 67.100 ;
        RECT 99.000 67.100 99.400 67.200 ;
        RECT 99.800 67.100 100.200 67.200 ;
        RECT 99.000 66.800 100.200 67.100 ;
        RECT 123.000 66.800 123.400 67.200 ;
        RECT 126.200 67.100 126.600 67.200 ;
        RECT 128.600 67.100 129.000 67.200 ;
        RECT 126.200 66.800 129.000 67.100 ;
        RECT 129.400 67.100 129.800 67.200 ;
        RECT 136.600 67.100 137.000 67.200 ;
        RECT 129.400 66.800 137.000 67.100 ;
        RECT 144.600 67.100 145.000 67.200 ;
        RECT 149.400 67.100 149.800 67.200 ;
        RECT 150.200 67.100 150.600 67.200 ;
        RECT 144.600 66.800 150.600 67.100 ;
        RECT 151.800 67.100 152.200 67.200 ;
        RECT 152.600 67.100 153.000 67.200 ;
        RECT 151.800 66.800 153.000 67.100 ;
        RECT 153.400 67.100 153.800 67.200 ;
        RECT 158.200 67.100 158.600 67.200 ;
        RECT 153.400 66.800 158.600 67.100 ;
        RECT 165.400 66.800 165.800 67.200 ;
        RECT 166.200 67.100 166.600 67.200 ;
        RECT 169.400 67.100 169.800 67.200 ;
        RECT 166.200 66.800 169.800 67.100 ;
        RECT 186.200 67.100 186.600 67.200 ;
        RECT 191.000 67.100 191.400 67.200 ;
        RECT 196.600 67.100 197.000 67.200 ;
        RECT 203.000 67.100 203.400 67.200 ;
        RECT 186.200 66.800 203.400 67.100 ;
        RECT 5.400 66.100 5.800 66.200 ;
        RECT 11.800 66.100 12.200 66.200 ;
        RECT 5.400 65.800 12.200 66.100 ;
        RECT 13.400 66.100 13.800 66.200 ;
        RECT 14.200 66.100 14.600 66.200 ;
        RECT 15.000 66.100 15.400 66.200 ;
        RECT 13.400 65.800 15.400 66.100 ;
        RECT 18.200 66.100 18.600 66.200 ;
        RECT 25.400 66.100 25.800 66.200 ;
        RECT 18.200 65.800 25.800 66.100 ;
        RECT 28.600 66.100 29.000 66.200 ;
        RECT 30.200 66.100 30.600 66.200 ;
        RECT 28.600 65.800 30.600 66.100 ;
        RECT 32.600 66.100 33.000 66.200 ;
        RECT 37.400 66.100 37.800 66.200 ;
        RECT 32.600 65.800 37.800 66.100 ;
        RECT 46.200 66.100 46.600 66.200 ;
        RECT 54.200 66.100 54.600 66.200 ;
        RECT 46.200 65.800 54.600 66.100 ;
        RECT 56.600 65.800 57.000 66.200 ;
        RECT 70.200 66.100 70.600 66.200 ;
        RECT 71.000 66.100 71.400 66.200 ;
        RECT 70.200 65.800 71.400 66.100 ;
        RECT 81.400 66.100 81.800 66.200 ;
        RECT 90.200 66.100 90.600 66.200 ;
        RECT 81.400 65.800 90.600 66.100 ;
        RECT 93.400 66.100 93.800 66.200 ;
        RECT 102.200 66.100 102.600 66.200 ;
        RECT 93.400 65.800 102.600 66.100 ;
        RECT 111.000 66.100 111.400 66.200 ;
        RECT 131.000 66.100 131.400 66.200 ;
        RECT 111.000 65.800 131.400 66.100 ;
        RECT 132.600 66.100 133.000 66.200 ;
        RECT 135.800 66.100 136.200 66.200 ;
        RECT 132.600 65.800 136.200 66.100 ;
        RECT 137.400 66.100 137.800 66.200 ;
        RECT 151.000 66.100 151.400 66.200 ;
        RECT 161.400 66.100 161.800 66.200 ;
        RECT 137.400 65.800 161.800 66.100 ;
        RECT 164.600 66.100 165.000 66.200 ;
        RECT 165.400 66.100 165.700 66.800 ;
        RECT 164.600 65.800 165.700 66.100 ;
        RECT 167.800 66.100 168.200 66.200 ;
        RECT 168.600 66.100 169.000 66.200 ;
        RECT 167.800 65.800 169.000 66.100 ;
        RECT 173.400 66.100 173.800 66.200 ;
        RECT 182.200 66.100 182.600 66.200 ;
        RECT 195.000 66.100 195.400 66.200 ;
        RECT 195.800 66.100 196.200 66.200 ;
        RECT 173.400 65.800 192.100 66.100 ;
        RECT 195.000 65.800 196.200 66.100 ;
        RECT 201.400 66.100 201.800 66.200 ;
        RECT 202.200 66.100 202.600 66.200 ;
        RECT 201.400 65.800 202.600 66.100 ;
        RECT 56.600 65.200 56.900 65.800 ;
        RECT 191.800 65.200 192.100 65.800 ;
        RECT 6.200 65.100 6.600 65.200 ;
        RECT 16.600 65.100 17.000 65.200 ;
        RECT 6.200 64.800 17.000 65.100 ;
        RECT 28.600 65.100 29.000 65.200 ;
        RECT 32.600 65.100 33.000 65.200 ;
        RECT 28.600 64.800 33.000 65.100 ;
        RECT 52.600 64.800 53.000 65.200 ;
        RECT 55.000 65.100 55.400 65.200 ;
        RECT 55.800 65.100 56.200 65.200 ;
        RECT 55.000 64.800 56.200 65.100 ;
        RECT 56.600 64.800 57.000 65.200 ;
        RECT 73.400 65.100 73.800 65.200 ;
        RECT 83.800 65.100 84.200 65.200 ;
        RECT 73.400 64.800 84.200 65.100 ;
        RECT 95.800 65.100 96.200 65.200 ;
        RECT 96.600 65.100 97.000 65.200 ;
        RECT 95.800 64.800 97.000 65.100 ;
        RECT 104.600 65.100 105.000 65.200 ;
        RECT 112.600 65.100 113.000 65.200 ;
        RECT 124.600 65.100 125.000 65.200 ;
        RECT 104.600 64.800 125.000 65.100 ;
        RECT 127.000 65.100 127.400 65.200 ;
        RECT 131.800 65.100 132.200 65.200 ;
        RECT 133.400 65.100 133.800 65.200 ;
        RECT 137.400 65.100 137.800 65.200 ;
        RECT 127.000 64.800 137.800 65.100 ;
        RECT 147.800 65.100 148.200 65.200 ;
        RECT 163.800 65.100 164.200 65.200 ;
        RECT 147.800 64.800 164.200 65.100 ;
        RECT 168.600 65.100 169.000 65.200 ;
        RECT 175.800 65.100 176.200 65.200 ;
        RECT 168.600 64.800 176.200 65.100 ;
        RECT 177.400 65.100 177.800 65.200 ;
        RECT 188.600 65.100 189.000 65.200 ;
        RECT 177.400 64.800 189.000 65.100 ;
        RECT 191.800 64.800 192.200 65.200 ;
        RECT 31.000 64.100 31.400 64.200 ;
        RECT 32.600 64.100 33.000 64.200 ;
        RECT 42.200 64.100 42.600 64.200 ;
        RECT 46.200 64.100 46.600 64.200 ;
        RECT 31.000 63.800 33.000 64.100 ;
        RECT 41.400 63.800 46.600 64.100 ;
        RECT 52.600 64.100 52.900 64.800 ;
        RECT 58.200 64.100 58.600 64.200 ;
        RECT 84.600 64.100 85.000 64.200 ;
        RECT 52.600 63.800 58.600 64.100 ;
        RECT 77.400 63.800 85.000 64.100 ;
        RECT 86.200 64.100 86.600 64.200 ;
        RECT 88.600 64.100 89.000 64.200 ;
        RECT 86.200 63.800 89.000 64.100 ;
        RECT 93.400 64.100 93.800 64.200 ;
        RECT 163.000 64.100 163.400 64.200 ;
        RECT 93.400 63.800 163.400 64.100 ;
        RECT 165.400 64.100 165.800 64.200 ;
        RECT 175.000 64.100 175.400 64.200 ;
        RECT 165.400 63.800 175.400 64.100 ;
        RECT 184.600 64.100 185.000 64.200 ;
        RECT 191.000 64.100 191.400 64.200 ;
        RECT 184.600 63.800 191.400 64.100 ;
        RECT 77.400 63.200 77.700 63.800 ;
        RECT 41.400 63.100 41.800 63.200 ;
        RECT 74.200 63.100 74.600 63.200 ;
        RECT 41.400 62.800 74.600 63.100 ;
        RECT 77.400 62.800 77.800 63.200 ;
        RECT 85.400 63.100 85.800 63.200 ;
        RECT 103.800 63.100 104.200 63.200 ;
        RECT 85.400 62.800 104.200 63.100 ;
        RECT 123.800 63.100 124.200 63.200 ;
        RECT 192.600 63.100 193.000 63.200 ;
        RECT 123.800 62.800 193.000 63.100 ;
        RECT 30.200 62.100 30.600 62.200 ;
        RECT 66.200 62.100 66.600 62.200 ;
        RECT 83.800 62.100 84.200 62.200 ;
        RECT 30.200 61.800 64.900 62.100 ;
        RECT 66.200 61.800 84.200 62.100 ;
        RECT 87.800 62.100 88.200 62.200 ;
        RECT 90.200 62.100 90.600 62.200 ;
        RECT 87.800 61.800 90.600 62.100 ;
        RECT 107.000 62.100 107.400 62.200 ;
        RECT 126.200 62.100 126.600 62.200 ;
        RECT 107.000 61.800 126.600 62.100 ;
        RECT 127.800 62.100 128.200 62.200 ;
        RECT 135.000 62.100 135.400 62.200 ;
        RECT 127.800 61.800 135.400 62.100 ;
        RECT 135.800 62.100 136.200 62.200 ;
        RECT 176.600 62.100 177.000 62.200 ;
        RECT 135.800 61.800 177.000 62.100 ;
        RECT 189.400 62.100 189.800 62.200 ;
        RECT 195.000 62.100 195.400 62.200 ;
        RECT 189.400 61.800 195.400 62.100 ;
        RECT 9.400 61.100 9.800 61.200 ;
        RECT 44.600 61.100 45.000 61.200 ;
        RECT 9.400 60.800 45.000 61.100 ;
        RECT 59.800 61.100 60.200 61.200 ;
        RECT 62.200 61.100 62.600 61.200 ;
        RECT 59.800 60.800 62.600 61.100 ;
        RECT 64.600 61.100 64.900 61.800 ;
        RECT 88.600 61.100 89.000 61.200 ;
        RECT 115.000 61.100 115.400 61.200 ;
        RECT 139.000 61.100 139.400 61.200 ;
        RECT 64.600 60.800 139.400 61.100 ;
        RECT 79.000 60.100 79.400 60.200 ;
        RECT 87.000 60.100 87.400 60.200 ;
        RECT 79.000 59.800 87.400 60.100 ;
        RECT 98.200 60.100 98.600 60.200 ;
        RECT 141.400 60.100 141.800 60.200 ;
        RECT 98.200 59.800 141.800 60.100 ;
        RECT 12.600 59.100 13.000 59.200 ;
        RECT 26.200 59.100 26.600 59.200 ;
        RECT 38.200 59.100 38.600 59.200 ;
        RECT 12.600 58.800 38.600 59.100 ;
        RECT 43.000 59.100 43.400 59.200 ;
        RECT 60.600 59.100 61.000 59.200 ;
        RECT 68.600 59.100 69.000 59.200 ;
        RECT 43.000 58.800 69.000 59.100 ;
        RECT 103.800 59.100 104.200 59.200 ;
        RECT 118.200 59.100 118.600 59.200 ;
        RECT 136.600 59.100 137.000 59.200 ;
        RECT 148.600 59.100 149.000 59.200 ;
        RECT 103.800 58.800 149.000 59.100 ;
        RECT 153.400 59.100 153.800 59.200 ;
        RECT 167.000 59.100 167.400 59.200 ;
        RECT 153.400 58.800 167.400 59.100 ;
        RECT 24.600 58.100 25.000 58.200 ;
        RECT 41.400 58.100 41.800 58.200 ;
        RECT 24.600 57.800 41.800 58.100 ;
        RECT 47.000 58.100 47.400 58.200 ;
        RECT 57.400 58.100 57.800 58.200 ;
        RECT 63.000 58.100 63.400 58.200 ;
        RECT 47.000 57.800 63.400 58.100 ;
        RECT 76.600 58.100 77.000 58.200 ;
        RECT 79.000 58.100 79.400 58.200 ;
        RECT 81.400 58.100 81.800 58.200 ;
        RECT 76.600 57.800 81.800 58.100 ;
        RECT 101.400 58.100 101.800 58.200 ;
        RECT 116.600 58.100 117.000 58.200 ;
        RECT 101.400 57.800 117.000 58.100 ;
        RECT 116.600 57.200 116.900 57.800 ;
        RECT 14.200 57.100 14.600 57.200 ;
        RECT 21.400 57.100 21.800 57.200 ;
        RECT 14.200 56.800 21.800 57.100 ;
        RECT 34.200 57.100 34.600 57.200 ;
        RECT 35.000 57.100 35.400 57.200 ;
        RECT 34.200 56.800 35.400 57.100 ;
        RECT 47.000 57.100 47.400 57.200 ;
        RECT 56.600 57.100 57.000 57.200 ;
        RECT 47.000 56.800 57.000 57.100 ;
        RECT 58.200 56.800 58.600 57.200 ;
        RECT 63.000 57.100 63.400 57.200 ;
        RECT 83.000 57.100 83.400 57.200 ;
        RECT 84.600 57.100 85.000 57.200 ;
        RECT 63.000 56.800 85.000 57.100 ;
        RECT 103.000 57.100 103.400 57.200 ;
        RECT 110.200 57.100 110.600 57.200 ;
        RECT 103.000 56.800 110.600 57.100 ;
        RECT 116.600 56.800 117.000 57.200 ;
        RECT 200.600 56.800 201.000 57.200 ;
        RECT 58.200 56.200 58.500 56.800 ;
        RECT 200.600 56.200 200.900 56.800 ;
        RECT 18.200 56.100 18.600 56.200 ;
        RECT 19.800 56.100 20.200 56.200 ;
        RECT 22.200 56.100 22.600 56.200 ;
        RECT 18.200 55.800 22.600 56.100 ;
        RECT 34.200 56.100 34.600 56.200 ;
        RECT 37.400 56.100 37.800 56.200 ;
        RECT 39.800 56.100 40.200 56.200 ;
        RECT 34.200 55.800 40.200 56.100 ;
        RECT 40.600 56.100 41.000 56.200 ;
        RECT 51.000 56.100 51.400 56.200 ;
        RECT 40.600 55.800 51.400 56.100 ;
        RECT 55.800 56.100 56.200 56.200 ;
        RECT 58.200 56.100 58.600 56.200 ;
        RECT 87.800 56.100 88.200 56.200 ;
        RECT 89.400 56.100 89.800 56.200 ;
        RECT 91.000 56.100 91.400 56.200 ;
        RECT 55.800 55.800 91.400 56.100 ;
        RECT 92.600 56.100 93.000 56.200 ;
        RECT 96.600 56.100 97.000 56.200 ;
        RECT 92.600 55.800 97.000 56.100 ;
        RECT 110.200 56.100 110.600 56.200 ;
        RECT 119.000 56.100 119.400 56.200 ;
        RECT 110.200 55.800 119.400 56.100 ;
        RECT 130.200 56.100 130.600 56.200 ;
        RECT 136.600 56.100 137.000 56.200 ;
        RECT 130.200 55.800 137.000 56.100 ;
        RECT 164.600 56.100 165.000 56.200 ;
        RECT 169.400 56.100 169.800 56.200 ;
        RECT 164.600 55.800 169.800 56.100 ;
        RECT 192.600 56.100 193.000 56.200 ;
        RECT 200.600 56.100 201.000 56.200 ;
        RECT 192.600 55.800 201.000 56.100 ;
        RECT 19.000 55.100 19.400 55.200 ;
        RECT 24.600 55.100 25.000 55.200 ;
        RECT 19.000 54.800 25.000 55.100 ;
        RECT 30.200 55.100 30.600 55.200 ;
        RECT 37.400 55.100 37.800 55.200 ;
        RECT 30.200 54.800 37.800 55.100 ;
        RECT 52.600 55.100 53.000 55.200 ;
        RECT 59.000 55.100 59.400 55.200 ;
        RECT 59.800 55.100 60.200 55.200 ;
        RECT 71.000 55.100 71.400 55.200 ;
        RECT 76.600 55.100 77.000 55.200 ;
        RECT 52.600 54.800 60.200 55.100 ;
        RECT 62.200 54.800 65.700 55.100 ;
        RECT 71.000 54.800 77.000 55.100 ;
        RECT 77.400 55.100 77.800 55.200 ;
        RECT 79.800 55.100 80.200 55.200 ;
        RECT 111.800 55.100 112.200 55.200 ;
        RECT 113.400 55.100 113.800 55.200 ;
        RECT 77.400 54.800 113.800 55.100 ;
        RECT 116.600 55.100 117.000 55.200 ;
        RECT 119.000 55.100 119.400 55.200 ;
        RECT 129.400 55.100 129.800 55.200 ;
        RECT 116.600 54.800 129.800 55.100 ;
        RECT 133.400 54.800 133.800 55.200 ;
        RECT 139.800 55.100 140.200 55.200 ;
        RECT 151.000 55.100 151.400 55.200 ;
        RECT 139.800 54.800 151.400 55.100 ;
        RECT 159.000 55.100 159.400 55.200 ;
        RECT 174.200 55.100 174.600 55.200 ;
        RECT 179.800 55.100 180.200 55.200 ;
        RECT 186.200 55.100 186.600 55.200 ;
        RECT 159.000 54.800 170.500 55.100 ;
        RECT 174.200 54.800 186.600 55.100 ;
        RECT 188.600 55.100 189.000 55.200 ;
        RECT 190.200 55.100 190.600 55.200 ;
        RECT 192.600 55.100 193.000 55.200 ;
        RECT 188.600 54.800 193.000 55.100 ;
        RECT 194.200 55.100 194.600 55.200 ;
        RECT 196.600 55.100 197.000 55.200 ;
        RECT 203.800 55.100 204.200 55.200 ;
        RECT 194.200 54.800 204.200 55.100 ;
        RECT 62.200 54.200 62.500 54.800 ;
        RECT 65.400 54.200 65.700 54.800 ;
        RECT 3.000 54.100 3.400 54.200 ;
        RECT 13.400 54.100 13.800 54.200 ;
        RECT 19.800 54.100 20.200 54.200 ;
        RECT 3.000 53.800 11.300 54.100 ;
        RECT 13.400 53.800 20.200 54.100 ;
        RECT 39.000 54.100 39.400 54.200 ;
        RECT 59.800 54.100 60.200 54.200 ;
        RECT 39.000 53.800 60.200 54.100 ;
        RECT 62.200 53.800 62.600 54.200 ;
        RECT 63.000 54.100 63.400 54.200 ;
        RECT 63.800 54.100 64.200 54.200 ;
        RECT 63.000 53.800 64.200 54.100 ;
        RECT 65.400 53.800 65.800 54.200 ;
        RECT 75.000 54.100 75.400 54.200 ;
        RECT 111.800 54.100 112.200 54.200 ;
        RECT 115.800 54.100 116.200 54.200 ;
        RECT 75.000 53.800 116.200 54.100 ;
        RECT 117.400 54.100 117.800 54.200 ;
        RECT 123.800 54.100 124.200 54.200 ;
        RECT 117.400 53.800 124.200 54.100 ;
        RECT 129.400 54.100 129.800 54.200 ;
        RECT 131.800 54.100 132.200 54.200 ;
        RECT 129.400 53.800 132.200 54.100 ;
        RECT 133.400 54.100 133.700 54.800 ;
        RECT 170.200 54.200 170.500 54.800 ;
        RECT 139.000 54.100 139.400 54.200 ;
        RECT 142.200 54.100 142.600 54.200 ;
        RECT 133.400 53.800 142.600 54.100 ;
        RECT 170.200 53.800 170.600 54.200 ;
        RECT 179.000 54.100 179.400 54.200 ;
        RECT 184.600 54.100 185.000 54.200 ;
        RECT 179.000 53.800 185.000 54.100 ;
        RECT 11.000 53.200 11.300 53.800 ;
        RECT 11.000 52.800 11.400 53.200 ;
        RECT 56.600 53.100 57.000 53.200 ;
        RECT 67.800 53.100 68.200 53.200 ;
        RECT 56.600 52.800 68.200 53.100 ;
        RECT 70.200 53.100 70.600 53.200 ;
        RECT 76.600 53.100 77.000 53.200 ;
        RECT 87.000 53.100 87.400 53.200 ;
        RECT 70.200 52.800 77.000 53.100 ;
        RECT 83.000 52.800 87.400 53.100 ;
        RECT 87.800 53.100 88.200 53.200 ;
        RECT 90.200 53.100 90.600 53.200 ;
        RECT 87.800 52.800 90.600 53.100 ;
        RECT 93.400 53.100 93.800 53.200 ;
        RECT 99.800 53.100 100.200 53.200 ;
        RECT 103.000 53.100 103.400 53.200 ;
        RECT 93.400 52.800 103.400 53.100 ;
        RECT 103.800 53.100 104.200 53.200 ;
        RECT 107.800 53.100 108.200 53.200 ;
        RECT 103.800 52.800 108.200 53.100 ;
        RECT 112.600 52.800 113.000 53.200 ;
        RECT 116.600 53.100 117.000 53.200 ;
        RECT 117.400 53.100 117.800 53.200 ;
        RECT 116.600 52.800 117.800 53.100 ;
        RECT 133.400 53.100 133.800 53.200 ;
        RECT 143.800 53.100 144.200 53.200 ;
        RECT 163.800 53.100 164.200 53.200 ;
        RECT 133.400 52.800 164.200 53.100 ;
        RECT 166.200 53.100 166.600 53.200 ;
        RECT 171.000 53.100 171.400 53.200 ;
        RECT 166.200 52.800 171.400 53.100 ;
        RECT 175.000 53.100 175.400 53.200 ;
        RECT 199.000 53.100 199.400 53.200 ;
        RECT 175.000 52.800 199.400 53.100 ;
        RECT 202.200 53.100 202.600 53.200 ;
        RECT 203.000 53.100 203.400 53.200 ;
        RECT 202.200 52.800 203.400 53.100 ;
        RECT 83.000 52.200 83.300 52.800 ;
        RECT 7.800 52.100 8.200 52.200 ;
        RECT 8.600 52.100 9.000 52.200 ;
        RECT 7.800 51.800 9.000 52.100 ;
        RECT 83.000 51.800 83.400 52.200 ;
        RECT 83.800 52.100 84.200 52.200 ;
        RECT 104.600 52.100 105.000 52.200 ;
        RECT 83.800 51.800 105.000 52.100 ;
        RECT 105.400 52.100 105.800 52.200 ;
        RECT 110.200 52.100 110.600 52.200 ;
        RECT 105.400 51.800 110.600 52.100 ;
        RECT 112.600 52.100 112.900 52.800 ;
        RECT 117.400 52.100 117.800 52.200 ;
        RECT 112.600 51.800 117.800 52.100 ;
        RECT 129.400 52.100 129.800 52.200 ;
        RECT 159.000 52.100 159.400 52.200 ;
        RECT 129.400 51.800 159.400 52.100 ;
        RECT 3.800 51.100 4.200 51.200 ;
        RECT 11.000 51.100 11.400 51.200 ;
        RECT 3.800 50.800 11.400 51.100 ;
        RECT 12.600 51.100 13.000 51.200 ;
        RECT 39.000 51.100 39.400 51.200 ;
        RECT 12.600 50.800 39.400 51.100 ;
        RECT 57.400 51.100 57.800 51.200 ;
        RECT 59.000 51.100 59.400 51.200 ;
        RECT 57.400 50.800 59.400 51.100 ;
        RECT 59.800 51.100 60.200 51.200 ;
        RECT 83.800 51.100 84.200 51.200 ;
        RECT 59.800 50.800 84.200 51.100 ;
        RECT 84.600 51.100 85.000 51.200 ;
        RECT 88.600 51.100 89.000 51.200 ;
        RECT 91.800 51.100 92.200 51.200 ;
        RECT 84.600 50.800 92.200 51.100 ;
        RECT 108.600 50.800 109.000 51.200 ;
        RECT 114.200 51.100 114.600 51.200 ;
        RECT 115.000 51.100 115.400 51.200 ;
        RECT 114.200 50.800 115.400 51.100 ;
        RECT 117.400 51.100 117.800 51.200 ;
        RECT 122.200 51.100 122.600 51.200 ;
        RECT 117.400 50.800 122.600 51.100 ;
        RECT 132.600 51.100 133.000 51.200 ;
        RECT 159.800 51.100 160.200 51.200 ;
        RECT 132.600 50.800 160.200 51.100 ;
        RECT 167.000 51.100 167.400 51.200 ;
        RECT 174.200 51.100 174.600 51.200 ;
        RECT 167.000 50.800 174.600 51.100 ;
        RECT 108.600 50.200 108.900 50.800 ;
        RECT 72.600 50.100 73.000 50.200 ;
        RECT 87.000 50.100 87.400 50.200 ;
        RECT 72.600 49.800 87.400 50.100 ;
        RECT 90.200 50.100 90.600 50.200 ;
        RECT 95.800 50.100 96.200 50.200 ;
        RECT 90.200 49.800 96.200 50.100 ;
        RECT 104.600 50.100 105.000 50.200 ;
        RECT 107.800 50.100 108.200 50.200 ;
        RECT 104.600 49.800 108.200 50.100 ;
        RECT 108.600 49.800 109.000 50.200 ;
        RECT 111.000 50.100 111.400 50.200 ;
        RECT 117.400 50.100 117.800 50.200 ;
        RECT 111.000 49.800 117.800 50.100 ;
        RECT 170.200 50.100 170.600 50.200 ;
        RECT 191.800 50.100 192.200 50.200 ;
        RECT 170.200 49.800 192.200 50.100 ;
        RECT 192.600 50.100 193.000 50.200 ;
        RECT 201.400 50.100 201.800 50.200 ;
        RECT 192.600 49.800 201.800 50.100 ;
        RECT 23.800 49.100 24.200 49.200 ;
        RECT 32.600 49.100 33.000 49.200 ;
        RECT 51.800 49.100 52.200 49.200 ;
        RECT 23.800 48.800 52.200 49.100 ;
        RECT 53.400 49.100 53.800 49.200 ;
        RECT 60.600 49.100 61.000 49.200 ;
        RECT 53.400 48.800 61.000 49.100 ;
        RECT 87.000 49.100 87.400 49.200 ;
        RECT 87.800 49.100 88.200 49.200 ;
        RECT 87.000 48.800 88.200 49.100 ;
        RECT 91.000 49.100 91.400 49.200 ;
        RECT 91.800 49.100 92.200 49.200 ;
        RECT 95.000 49.100 95.400 49.200 ;
        RECT 109.400 49.100 109.800 49.200 ;
        RECT 91.000 48.800 92.200 49.100 ;
        RECT 94.200 48.800 109.800 49.100 ;
        RECT 114.200 49.100 114.600 49.200 ;
        RECT 135.000 49.100 135.400 49.200 ;
        RECT 143.800 49.100 144.200 49.200 ;
        RECT 114.200 48.800 144.200 49.100 ;
        RECT 145.400 49.100 145.800 49.200 ;
        RECT 151.800 49.100 152.200 49.200 ;
        RECT 161.400 49.100 161.800 49.200 ;
        RECT 167.000 49.100 167.400 49.200 ;
        RECT 145.400 48.800 167.400 49.100 ;
        RECT 22.200 48.100 22.600 48.200 ;
        RECT 31.800 48.100 32.200 48.200 ;
        RECT 35.000 48.100 35.400 48.200 ;
        RECT 22.200 47.800 35.400 48.100 ;
        RECT 39.000 48.100 39.400 48.200 ;
        RECT 64.600 48.100 65.000 48.200 ;
        RECT 39.000 47.800 65.000 48.100 ;
        RECT 75.000 48.100 75.400 48.200 ;
        RECT 82.200 48.100 82.600 48.200 ;
        RECT 75.000 47.800 82.600 48.100 ;
        RECT 83.000 48.100 83.400 48.200 ;
        RECT 133.400 48.100 133.800 48.200 ;
        RECT 83.000 47.800 133.800 48.100 ;
        RECT 147.800 47.800 148.200 48.200 ;
        RECT 148.600 48.100 149.000 48.200 ;
        RECT 150.200 48.100 150.600 48.200 ;
        RECT 148.600 47.800 150.600 48.100 ;
        RECT 178.200 48.100 178.600 48.200 ;
        RECT 188.600 48.100 189.000 48.200 ;
        RECT 178.200 47.800 189.000 48.100 ;
        RECT 195.000 48.100 195.400 48.200 ;
        RECT 201.400 48.100 201.800 48.200 ;
        RECT 202.200 48.100 202.600 48.200 ;
        RECT 195.000 47.800 202.600 48.100 ;
        RECT 45.400 47.200 45.700 47.800 ;
        RECT 147.800 47.200 148.100 47.800 ;
        RECT 9.400 47.100 9.800 47.200 ;
        RECT 12.600 47.100 13.000 47.200 ;
        RECT 9.400 46.800 13.000 47.100 ;
        RECT 37.400 47.100 37.800 47.200 ;
        RECT 42.200 47.100 42.600 47.200 ;
        RECT 37.400 46.800 42.600 47.100 ;
        RECT 45.400 46.800 45.800 47.200 ;
        RECT 49.400 47.100 49.800 47.200 ;
        RECT 77.400 47.100 77.800 47.200 ;
        RECT 49.400 46.800 77.800 47.100 ;
        RECT 80.600 46.800 81.000 47.200 ;
        RECT 84.600 47.100 85.000 47.200 ;
        RECT 92.600 47.100 93.000 47.200 ;
        RECT 84.600 46.800 93.000 47.100 ;
        RECT 95.000 47.100 95.400 47.200 ;
        RECT 103.800 47.100 104.200 47.200 ;
        RECT 95.000 46.800 104.200 47.100 ;
        RECT 104.600 47.100 105.000 47.200 ;
        RECT 105.400 47.100 105.800 47.200 ;
        RECT 104.600 46.800 105.800 47.100 ;
        RECT 106.200 47.100 106.600 47.200 ;
        RECT 107.800 47.100 108.200 47.200 ;
        RECT 106.200 46.800 108.200 47.100 ;
        RECT 108.600 47.100 109.000 47.200 ;
        RECT 112.600 47.100 113.000 47.200 ;
        RECT 108.600 46.800 113.000 47.100 ;
        RECT 113.400 47.100 113.800 47.200 ;
        RECT 127.800 47.100 128.200 47.200 ;
        RECT 113.400 46.800 128.200 47.100 ;
        RECT 140.600 46.800 141.000 47.200 ;
        RECT 145.400 47.100 145.800 47.200 ;
        RECT 147.800 47.100 148.200 47.200 ;
        RECT 145.400 46.800 148.200 47.100 ;
        RECT 148.600 47.100 149.000 47.200 ;
        RECT 155.000 47.100 155.400 47.200 ;
        RECT 148.600 46.800 155.400 47.100 ;
        RECT 159.800 47.100 160.200 47.200 ;
        RECT 190.200 47.100 190.600 47.200 ;
        RECT 159.800 46.800 190.600 47.100 ;
        RECT 202.200 47.100 202.600 47.200 ;
        RECT 203.000 47.100 203.400 47.200 ;
        RECT 202.200 46.800 203.400 47.100 ;
        RECT 11.800 46.100 12.200 46.200 ;
        RECT 12.600 46.100 13.000 46.200 ;
        RECT 11.800 45.800 13.000 46.100 ;
        RECT 15.000 46.100 15.400 46.200 ;
        RECT 16.600 46.100 17.000 46.200 ;
        RECT 15.000 45.800 17.000 46.100 ;
        RECT 22.200 46.100 22.600 46.200 ;
        RECT 27.800 46.100 28.200 46.300 ;
        RECT 22.200 45.900 28.200 46.100 ;
        RECT 35.000 46.100 35.400 46.200 ;
        RECT 37.400 46.100 37.800 46.200 ;
        RECT 22.200 45.800 28.100 45.900 ;
        RECT 35.000 45.800 37.800 46.100 ;
        RECT 44.600 46.100 45.000 46.200 ;
        RECT 61.400 46.100 61.800 46.200 ;
        RECT 71.000 46.100 71.400 46.200 ;
        RECT 44.600 45.800 71.400 46.100 ;
        RECT 80.600 46.100 80.900 46.800 ;
        RECT 84.600 46.100 84.900 46.800 ;
        RECT 80.600 45.800 84.900 46.100 ;
        RECT 86.200 45.800 86.600 46.200 ;
        RECT 95.800 46.100 96.200 46.200 ;
        RECT 96.600 46.100 97.000 46.200 ;
        RECT 95.800 45.800 97.000 46.100 ;
        RECT 97.400 46.100 97.800 46.200 ;
        RECT 98.200 46.100 98.600 46.200 ;
        RECT 97.400 45.800 98.600 46.100 ;
        RECT 100.600 46.100 101.000 46.200 ;
        RECT 105.400 46.100 105.800 46.200 ;
        RECT 100.600 45.800 105.800 46.100 ;
        RECT 107.000 46.100 107.400 46.200 ;
        RECT 112.600 46.100 113.000 46.200 ;
        RECT 116.600 46.100 117.000 46.200 ;
        RECT 130.200 46.100 130.600 46.200 ;
        RECT 138.200 46.100 138.600 46.200 ;
        RECT 107.000 45.800 138.600 46.100 ;
        RECT 140.600 46.100 140.900 46.800 ;
        RECT 146.200 46.100 146.600 46.200 ;
        RECT 140.600 45.800 146.600 46.100 ;
        RECT 149.400 46.100 149.800 46.200 ;
        RECT 164.600 46.100 165.000 46.200 ;
        RECT 177.400 46.100 177.800 46.200 ;
        RECT 149.400 45.800 177.800 46.100 ;
        RECT 184.600 46.100 185.000 46.200 ;
        RECT 187.800 46.100 188.200 46.200 ;
        RECT 184.600 45.800 188.200 46.100 ;
        RECT 195.800 46.100 196.200 46.200 ;
        RECT 200.600 46.100 201.000 46.200 ;
        RECT 195.800 45.800 201.000 46.100 ;
        RECT 201.400 46.100 201.800 46.200 ;
        RECT 203.800 46.100 204.200 46.200 ;
        RECT 201.400 45.800 204.200 46.100 ;
        RECT 86.200 45.200 86.500 45.800 ;
        RECT 18.200 45.100 18.600 45.200 ;
        RECT 23.000 45.100 23.400 45.200 ;
        RECT 49.400 45.100 49.800 45.200 ;
        RECT 18.200 44.800 49.800 45.100 ;
        RECT 52.600 45.100 53.000 45.200 ;
        RECT 55.000 45.100 55.400 45.200 ;
        RECT 82.200 45.100 82.600 45.200 ;
        RECT 52.600 44.800 82.600 45.100 ;
        RECT 86.200 44.800 86.600 45.200 ;
        RECT 89.400 45.100 89.800 45.200 ;
        RECT 93.400 45.100 93.800 45.200 ;
        RECT 89.400 44.800 93.800 45.100 ;
        RECT 99.800 45.100 100.200 45.200 ;
        RECT 103.000 45.100 103.400 45.200 ;
        RECT 99.800 44.800 103.400 45.100 ;
        RECT 113.400 45.100 113.800 45.200 ;
        RECT 114.200 45.100 114.600 45.200 ;
        RECT 115.800 45.100 116.200 45.200 ;
        RECT 113.400 44.800 116.200 45.100 ;
        RECT 126.200 45.100 126.600 45.200 ;
        RECT 127.000 45.100 127.400 45.200 ;
        RECT 126.200 44.800 127.400 45.100 ;
        RECT 127.800 44.800 128.200 45.200 ;
        RECT 148.600 45.100 149.000 45.200 ;
        RECT 149.400 45.100 149.800 45.200 ;
        RECT 148.600 44.800 149.800 45.100 ;
        RECT 155.800 45.100 156.200 45.200 ;
        RECT 164.600 45.100 165.000 45.200 ;
        RECT 155.800 44.800 165.000 45.100 ;
        RECT 127.800 44.200 128.100 44.800 ;
        RECT 19.000 44.100 19.400 44.200 ;
        RECT 22.200 44.100 22.600 44.200 ;
        RECT 19.000 43.800 22.600 44.100 ;
        RECT 51.800 44.100 52.200 44.200 ;
        RECT 53.400 44.100 53.800 44.200 ;
        RECT 51.800 43.800 53.800 44.100 ;
        RECT 75.000 44.100 75.400 44.200 ;
        RECT 98.200 44.100 98.600 44.200 ;
        RECT 75.000 43.800 98.600 44.100 ;
        RECT 103.800 44.100 104.200 44.200 ;
        RECT 108.600 44.100 109.000 44.200 ;
        RECT 103.800 43.800 109.000 44.100 ;
        RECT 127.800 43.800 128.200 44.200 ;
        RECT 151.000 44.100 151.400 44.200 ;
        RECT 156.600 44.100 157.000 44.200 ;
        RECT 151.000 43.800 157.000 44.100 ;
        RECT 162.200 44.100 162.600 44.200 ;
        RECT 164.600 44.100 165.000 44.200 ;
        RECT 162.200 43.800 165.000 44.100 ;
        RECT 43.800 43.100 44.200 43.200 ;
        RECT 56.600 43.100 57.000 43.200 ;
        RECT 43.800 42.800 57.000 43.100 ;
        RECT 69.400 43.100 69.800 43.200 ;
        RECT 89.400 43.100 89.800 43.200 ;
        RECT 69.400 42.800 89.800 43.100 ;
        RECT 90.200 43.100 90.600 43.200 ;
        RECT 105.400 43.100 105.800 43.200 ;
        RECT 122.200 43.100 122.600 43.200 ;
        RECT 90.200 42.800 122.600 43.100 ;
        RECT 148.600 43.100 149.000 43.200 ;
        RECT 165.400 43.100 165.800 43.200 ;
        RECT 191.800 43.100 192.200 43.200 ;
        RECT 148.600 42.800 192.200 43.100 ;
        RECT 40.600 42.100 41.000 42.200 ;
        RECT 43.800 42.100 44.200 42.200 ;
        RECT 40.600 41.800 44.200 42.100 ;
        RECT 51.000 42.100 51.400 42.200 ;
        RECT 63.000 42.100 63.400 42.200 ;
        RECT 51.000 41.800 63.400 42.100 ;
        RECT 84.600 42.100 85.000 42.200 ;
        RECT 165.400 42.100 165.800 42.200 ;
        RECT 167.800 42.100 168.200 42.200 ;
        RECT 84.600 41.800 168.200 42.100 ;
        RECT 170.200 42.100 170.600 42.200 ;
        RECT 171.000 42.100 171.400 42.200 ;
        RECT 170.200 41.800 171.400 42.100 ;
        RECT 174.200 42.100 174.600 42.200 ;
        RECT 184.600 42.100 185.000 42.200 ;
        RECT 174.200 41.800 185.000 42.100 ;
        RECT 186.200 42.100 186.600 42.200 ;
        RECT 187.000 42.100 187.400 42.200 ;
        RECT 186.200 41.800 187.400 42.100 ;
        RECT 190.200 42.100 190.600 42.200 ;
        RECT 191.800 42.100 192.200 42.200 ;
        RECT 190.200 41.800 192.200 42.100 ;
        RECT 64.600 41.100 65.000 41.200 ;
        RECT 75.000 41.100 75.400 41.200 ;
        RECT 64.600 40.800 75.400 41.100 ;
        RECT 82.200 41.100 82.600 41.200 ;
        RECT 119.000 41.100 119.400 41.200 ;
        RECT 82.200 40.800 119.400 41.100 ;
        RECT 155.000 41.100 155.400 41.200 ;
        RECT 173.400 41.100 173.800 41.200 ;
        RECT 155.000 40.800 173.800 41.100 ;
        RECT 57.400 40.100 57.800 40.200 ;
        RECT 62.200 40.100 62.600 40.200 ;
        RECT 73.400 40.100 73.800 40.200 ;
        RECT 83.000 40.100 83.400 40.200 ;
        RECT 57.400 39.800 83.400 40.100 ;
        RECT 89.400 40.100 89.800 40.200 ;
        RECT 106.200 40.100 106.600 40.200 ;
        RECT 89.400 39.800 106.600 40.100 ;
        RECT 109.400 40.100 109.800 40.200 ;
        RECT 111.000 40.100 111.400 40.200 ;
        RECT 109.400 39.800 111.400 40.100 ;
        RECT 124.600 40.100 125.000 40.200 ;
        RECT 139.800 40.100 140.200 40.200 ;
        RECT 124.600 39.800 140.200 40.100 ;
        RECT 162.200 40.100 162.600 40.200 ;
        RECT 167.800 40.100 168.200 40.200 ;
        RECT 162.200 39.800 168.200 40.100 ;
        RECT 11.800 39.100 12.200 39.200 ;
        RECT 13.400 39.100 13.800 39.200 ;
        RECT 38.200 39.100 38.600 39.200 ;
        RECT 11.800 38.800 38.600 39.100 ;
        RECT 68.600 39.100 69.000 39.200 ;
        RECT 84.600 39.100 85.000 39.200 ;
        RECT 87.000 39.100 87.400 39.200 ;
        RECT 128.600 39.100 129.000 39.200 ;
        RECT 68.600 38.800 129.000 39.100 ;
        RECT 132.600 39.100 133.000 39.200 ;
        RECT 154.200 39.100 154.600 39.200 ;
        RECT 132.600 38.800 154.600 39.100 ;
        RECT 160.600 39.100 161.000 39.200 ;
        RECT 163.000 39.100 163.400 39.200 ;
        RECT 160.600 38.800 163.400 39.100 ;
        RECT 167.000 39.100 167.400 39.200 ;
        RECT 195.800 39.100 196.200 39.200 ;
        RECT 167.000 38.800 196.200 39.100 ;
        RECT 31.800 38.100 32.200 38.200 ;
        RECT 51.800 38.100 52.200 38.200 ;
        RECT 31.800 37.800 52.200 38.100 ;
        RECT 61.400 38.100 61.800 38.200 ;
        RECT 159.000 38.100 159.400 38.200 ;
        RECT 162.200 38.100 162.600 38.200 ;
        RECT 61.400 37.800 135.300 38.100 ;
        RECT 159.000 37.800 162.600 38.100 ;
        RECT 169.400 38.100 169.800 38.200 ;
        RECT 171.800 38.100 172.200 38.200 ;
        RECT 169.400 37.800 181.700 38.100 ;
        RECT 5.400 37.100 5.800 37.200 ;
        RECT 15.800 37.100 16.200 37.200 ;
        RECT 5.400 36.800 16.200 37.100 ;
        RECT 19.800 37.100 20.200 37.200 ;
        RECT 28.600 37.100 29.000 37.200 ;
        RECT 19.800 36.800 29.000 37.100 ;
        RECT 31.800 37.100 32.100 37.800 ;
        RECT 135.000 37.200 135.300 37.800 ;
        RECT 181.400 37.200 181.700 37.800 ;
        RECT 35.800 37.100 36.200 37.200 ;
        RECT 31.800 36.800 36.200 37.100 ;
        RECT 37.400 36.800 37.800 37.200 ;
        RECT 39.800 36.800 40.200 37.200 ;
        RECT 75.000 36.800 75.400 37.200 ;
        RECT 80.600 36.800 81.000 37.200 ;
        RECT 82.200 37.100 82.600 37.200 ;
        RECT 85.400 37.100 85.800 37.200 ;
        RECT 98.200 37.100 98.600 37.200 ;
        RECT 82.200 36.800 98.600 37.100 ;
        RECT 99.000 37.100 99.400 37.200 ;
        RECT 100.600 37.100 101.000 37.200 ;
        RECT 99.000 36.800 101.000 37.100 ;
        RECT 108.600 37.100 109.000 37.200 ;
        RECT 109.400 37.100 109.800 37.200 ;
        RECT 111.800 37.100 112.200 37.200 ;
        RECT 108.600 36.800 109.800 37.100 ;
        RECT 110.200 36.800 112.200 37.100 ;
        RECT 113.400 37.100 113.800 37.200 ;
        RECT 120.600 37.100 121.000 37.200 ;
        RECT 113.400 36.800 121.000 37.100 ;
        RECT 135.000 37.100 135.400 37.200 ;
        RECT 136.600 37.100 137.000 37.200 ;
        RECT 135.000 36.800 137.000 37.100 ;
        RECT 164.600 37.100 165.000 37.200 ;
        RECT 173.400 37.100 173.800 37.200 ;
        RECT 164.600 36.800 173.800 37.100 ;
        RECT 181.400 37.100 181.800 37.200 ;
        RECT 183.800 37.100 184.200 37.200 ;
        RECT 194.200 37.100 194.600 37.200 ;
        RECT 181.400 36.800 194.600 37.100 ;
        RECT 37.400 36.200 37.700 36.800 ;
        RECT 39.800 36.200 40.100 36.800 ;
        RECT 75.000 36.200 75.300 36.800 ;
        RECT 80.600 36.200 80.900 36.800 ;
        RECT 15.800 36.100 16.200 36.200 ;
        RECT 16.600 36.100 17.000 36.200 ;
        RECT 15.800 35.800 17.000 36.100 ;
        RECT 18.200 35.800 18.600 36.200 ;
        RECT 28.600 36.100 29.000 36.200 ;
        RECT 32.600 36.100 33.000 36.200 ;
        RECT 37.400 36.100 37.800 36.200 ;
        RECT 28.600 35.800 37.800 36.100 ;
        RECT 39.800 36.100 40.200 36.200 ;
        RECT 43.000 36.100 43.400 36.200 ;
        RECT 39.800 35.800 43.400 36.100 ;
        RECT 46.200 36.100 46.600 36.200 ;
        RECT 47.800 36.100 48.200 36.200 ;
        RECT 46.200 35.800 48.200 36.100 ;
        RECT 55.800 36.100 56.200 36.200 ;
        RECT 59.800 36.100 60.200 36.200 ;
        RECT 63.800 36.100 64.200 36.200 ;
        RECT 55.800 35.800 64.200 36.100 ;
        RECT 64.600 35.800 65.000 36.200 ;
        RECT 65.400 36.100 65.800 36.200 ;
        RECT 67.000 36.100 67.400 36.200 ;
        RECT 65.400 35.800 67.400 36.100 ;
        RECT 75.000 35.800 75.400 36.200 ;
        RECT 80.600 36.100 81.000 36.200 ;
        RECT 110.200 36.100 110.500 36.800 ;
        RECT 80.600 35.800 110.500 36.100 ;
        RECT 135.800 36.100 136.200 36.200 ;
        RECT 155.800 36.100 156.200 36.200 ;
        RECT 135.800 35.800 156.200 36.100 ;
        RECT 156.600 36.100 157.000 36.200 ;
        RECT 174.200 36.100 174.600 36.200 ;
        RECT 178.200 36.100 178.600 36.200 ;
        RECT 189.400 36.100 189.800 36.200 ;
        RECT 156.600 35.800 178.600 36.100 ;
        RECT 179.000 35.800 189.800 36.100 ;
        RECT 18.200 35.200 18.500 35.800 ;
        RECT 64.600 35.200 64.900 35.800 ;
        RECT 1.400 35.100 1.800 35.200 ;
        RECT 14.200 35.100 14.600 35.200 ;
        RECT 17.400 35.100 17.800 35.200 ;
        RECT 1.400 34.800 17.800 35.100 ;
        RECT 18.200 34.800 18.600 35.200 ;
        RECT 27.800 35.100 28.200 35.200 ;
        RECT 35.000 35.100 35.400 35.200 ;
        RECT 27.800 34.800 35.400 35.100 ;
        RECT 39.800 35.100 40.200 35.200 ;
        RECT 40.600 35.100 41.000 35.200 ;
        RECT 39.800 34.800 41.000 35.100 ;
        RECT 64.600 34.800 65.000 35.200 ;
        RECT 65.400 35.100 65.800 35.200 ;
        RECT 70.200 35.100 70.600 35.200 ;
        RECT 65.400 34.800 70.600 35.100 ;
        RECT 71.000 35.100 71.400 35.200 ;
        RECT 77.400 35.100 77.800 35.200 ;
        RECT 95.000 35.100 95.400 35.200 ;
        RECT 71.000 34.800 95.400 35.100 ;
        RECT 97.400 34.800 97.800 35.200 ;
        RECT 98.200 35.100 98.600 35.200 ;
        RECT 111.000 35.100 111.400 35.200 ;
        RECT 98.200 34.800 111.400 35.100 ;
        RECT 128.600 35.100 129.000 35.200 ;
        RECT 130.200 35.100 130.600 35.200 ;
        RECT 169.400 35.100 169.800 35.200 ;
        RECT 128.600 34.800 169.800 35.100 ;
        RECT 177.400 35.100 177.800 35.200 ;
        RECT 179.000 35.100 179.300 35.800 ;
        RECT 177.400 34.800 179.300 35.100 ;
        RECT 180.600 35.100 181.000 35.200 ;
        RECT 180.600 34.800 188.900 35.100 ;
        RECT 17.400 34.100 17.800 34.200 ;
        RECT 19.000 34.100 19.400 34.200 ;
        RECT 29.400 34.100 29.800 34.200 ;
        RECT 17.400 33.800 29.800 34.100 ;
        RECT 30.200 34.100 30.600 34.200 ;
        RECT 43.800 34.100 44.200 34.200 ;
        RECT 30.200 33.800 44.200 34.100 ;
        RECT 48.600 34.100 49.000 34.200 ;
        RECT 49.400 34.100 49.800 34.200 ;
        RECT 48.600 33.800 49.800 34.100 ;
        RECT 53.400 34.100 53.800 34.200 ;
        RECT 58.200 34.100 58.600 34.200 ;
        RECT 53.400 33.800 58.600 34.100 ;
        RECT 61.400 34.100 61.800 34.200 ;
        RECT 66.200 34.100 66.600 34.200 ;
        RECT 68.600 34.100 69.000 34.200 ;
        RECT 61.400 33.800 69.000 34.100 ;
        RECT 71.800 34.100 72.200 34.200 ;
        RECT 83.800 34.100 84.200 34.200 ;
        RECT 71.800 33.800 84.200 34.100 ;
        RECT 87.000 34.100 87.400 34.200 ;
        RECT 93.400 34.100 93.800 34.200 ;
        RECT 87.000 33.800 93.800 34.100 ;
        RECT 97.400 34.100 97.700 34.800 ;
        RECT 188.600 34.200 188.900 34.800 ;
        RECT 99.800 34.100 100.200 34.200 ;
        RECT 97.400 33.800 100.200 34.100 ;
        RECT 105.400 34.100 105.800 34.200 ;
        RECT 106.200 34.100 106.600 34.200 ;
        RECT 105.400 33.800 106.600 34.100 ;
        RECT 110.200 34.100 110.600 34.200 ;
        RECT 113.400 34.100 113.800 34.200 ;
        RECT 115.000 34.100 115.400 34.200 ;
        RECT 110.200 33.800 115.400 34.100 ;
        RECT 120.600 34.100 121.000 34.200 ;
        RECT 127.800 34.100 128.200 34.200 ;
        RECT 120.600 33.800 128.200 34.100 ;
        RECT 133.400 34.100 133.800 34.200 ;
        RECT 142.200 34.100 142.600 34.200 ;
        RECT 169.400 34.100 169.800 34.200 ;
        RECT 133.400 33.800 142.600 34.100 ;
        RECT 166.200 33.800 169.800 34.100 ;
        RECT 179.000 33.800 179.400 34.200 ;
        RECT 188.600 33.800 189.000 34.200 ;
        RECT 166.200 33.200 166.500 33.800 ;
        RECT 10.200 33.100 10.600 33.200 ;
        RECT 15.800 33.100 16.200 33.200 ;
        RECT 10.200 32.800 16.200 33.100 ;
        RECT 39.000 32.800 39.400 33.200 ;
        RECT 43.800 33.100 44.200 33.200 ;
        RECT 46.200 33.100 46.600 33.200 ;
        RECT 57.400 33.100 57.800 33.200 ;
        RECT 71.000 33.100 71.400 33.200 ;
        RECT 43.800 32.800 71.400 33.100 ;
        RECT 75.800 33.100 76.200 33.200 ;
        RECT 79.800 33.100 80.200 33.200 ;
        RECT 99.000 33.100 99.400 33.200 ;
        RECT 115.800 33.100 116.200 33.200 ;
        RECT 75.800 32.800 116.200 33.100 ;
        RECT 116.600 33.100 117.000 33.200 ;
        RECT 143.000 33.100 143.400 33.200 ;
        RECT 116.600 32.800 143.400 33.100 ;
        RECT 166.200 32.800 166.600 33.200 ;
        RECT 179.000 33.100 179.300 33.800 ;
        RECT 184.600 33.100 185.000 33.200 ;
        RECT 179.000 32.800 185.000 33.100 ;
        RECT 197.400 33.100 197.800 33.200 ;
        RECT 201.400 33.100 201.800 33.200 ;
        RECT 197.400 32.800 201.800 33.100 ;
        RECT 7.000 32.100 7.400 32.200 ;
        RECT 12.600 32.100 13.000 32.200 ;
        RECT 7.000 31.800 13.000 32.100 ;
        RECT 16.600 32.100 17.000 32.200 ;
        RECT 19.800 32.100 20.200 32.200 ;
        RECT 16.600 31.800 20.200 32.100 ;
        RECT 29.400 32.100 29.800 32.200 ;
        RECT 33.400 32.100 33.800 32.200 ;
        RECT 29.400 31.800 33.800 32.100 ;
        RECT 39.000 32.100 39.300 32.800 ;
        RECT 47.000 32.100 47.400 32.200 ;
        RECT 39.000 31.800 47.400 32.100 ;
        RECT 69.400 32.100 69.800 32.200 ;
        RECT 77.400 32.100 77.800 32.200 ;
        RECT 69.400 31.800 77.800 32.100 ;
        RECT 78.200 32.100 78.600 32.200 ;
        RECT 80.600 32.100 81.000 32.200 ;
        RECT 78.200 31.800 81.000 32.100 ;
        RECT 82.200 32.100 82.600 32.200 ;
        RECT 99.000 32.100 99.400 32.200 ;
        RECT 82.200 31.800 99.400 32.100 ;
        RECT 100.600 32.100 101.000 32.200 ;
        RECT 103.800 32.100 104.200 32.200 ;
        RECT 100.600 31.800 104.200 32.100 ;
        RECT 104.600 32.100 105.000 32.200 ;
        RECT 105.400 32.100 105.800 32.200 ;
        RECT 104.600 31.800 105.800 32.100 ;
        RECT 106.200 32.100 106.600 32.200 ;
        RECT 112.600 32.100 113.000 32.200 ;
        RECT 106.200 31.800 113.000 32.100 ;
        RECT 130.200 32.100 130.600 32.200 ;
        RECT 136.600 32.100 137.000 32.200 ;
        RECT 130.200 31.800 137.000 32.100 ;
        RECT 172.600 32.100 173.000 32.200 ;
        RECT 176.600 32.100 177.000 32.200 ;
        RECT 181.400 32.100 181.800 32.200 ;
        RECT 172.600 31.800 181.800 32.100 ;
        RECT 28.600 31.100 29.000 31.200 ;
        RECT 54.200 31.100 54.600 31.200 ;
        RECT 28.600 30.800 54.600 31.100 ;
        RECT 59.000 31.100 59.400 31.200 ;
        RECT 96.600 31.100 97.000 31.200 ;
        RECT 59.000 30.800 97.000 31.100 ;
        RECT 111.800 31.100 112.200 31.200 ;
        RECT 142.200 31.100 142.600 31.200 ;
        RECT 161.400 31.100 161.800 31.200 ;
        RECT 111.800 30.800 161.800 31.100 ;
        RECT 196.600 31.100 197.000 31.200 ;
        RECT 197.400 31.100 197.800 31.200 ;
        RECT 196.600 30.800 197.800 31.100 ;
        RECT 41.400 30.100 41.800 30.200 ;
        RECT 50.200 30.100 50.600 30.200 ;
        RECT 41.400 29.800 50.600 30.100 ;
        RECT 51.000 30.100 51.400 30.200 ;
        RECT 55.000 30.100 55.400 30.200 ;
        RECT 61.400 30.100 61.800 30.200 ;
        RECT 67.000 30.100 67.400 30.200 ;
        RECT 71.800 30.100 72.200 30.200 ;
        RECT 77.400 30.100 77.800 30.200 ;
        RECT 83.000 30.100 83.400 30.200 ;
        RECT 51.000 29.800 83.400 30.100 ;
        RECT 115.000 30.100 115.400 30.200 ;
        RECT 119.000 30.100 119.400 30.200 ;
        RECT 115.000 29.800 119.400 30.100 ;
        RECT 151.000 30.100 151.400 30.200 ;
        RECT 157.400 30.100 157.800 30.200 ;
        RECT 151.000 29.800 157.800 30.100 ;
        RECT 179.800 30.100 180.200 30.200 ;
        RECT 187.000 30.100 187.400 30.200 ;
        RECT 179.800 29.800 187.400 30.100 ;
        RECT 31.000 29.100 31.400 29.200 ;
        RECT 34.200 29.100 34.600 29.200 ;
        RECT 35.000 29.100 35.400 29.200 ;
        RECT 31.000 28.800 35.400 29.100 ;
        RECT 46.200 29.100 46.600 29.200 ;
        RECT 82.200 29.100 82.600 29.200 ;
        RECT 107.800 29.100 108.200 29.200 ;
        RECT 171.000 29.100 171.400 29.200 ;
        RECT 46.200 28.800 171.400 29.100 ;
        RECT 171.800 29.100 172.200 29.200 ;
        RECT 179.000 29.100 179.400 29.200 ;
        RECT 171.800 28.800 179.400 29.100 ;
        RECT 23.000 28.100 23.400 28.200 ;
        RECT 32.600 28.100 33.000 28.200 ;
        RECT 23.000 27.800 33.000 28.100 ;
        RECT 35.800 27.800 36.200 28.200 ;
        RECT 43.800 28.100 44.200 28.200 ;
        RECT 49.400 28.100 49.800 28.200 ;
        RECT 63.000 28.100 63.400 28.200 ;
        RECT 81.400 28.100 81.800 28.200 ;
        RECT 43.800 27.800 61.700 28.100 ;
        RECT 63.000 27.800 81.800 28.100 ;
        RECT 83.000 27.800 83.400 28.200 ;
        RECT 85.400 28.100 85.800 28.200 ;
        RECT 87.000 28.100 87.400 28.200 ;
        RECT 85.400 27.800 87.400 28.100 ;
        RECT 87.800 28.100 88.200 28.200 ;
        RECT 93.400 28.100 93.800 28.200 ;
        RECT 87.800 27.800 93.800 28.100 ;
        RECT 95.000 27.800 95.400 28.200 ;
        RECT 104.600 27.800 105.000 28.200 ;
        RECT 111.800 27.800 112.200 28.200 ;
        RECT 117.400 27.800 117.800 28.200 ;
        RECT 121.400 28.100 121.800 28.200 ;
        RECT 144.600 28.100 145.000 28.200 ;
        RECT 159.800 28.100 160.200 28.200 ;
        RECT 121.400 27.800 160.200 28.100 ;
        RECT 163.000 28.100 163.400 28.200 ;
        RECT 167.000 28.100 167.400 28.200 ;
        RECT 163.000 27.800 167.400 28.100 ;
        RECT 167.800 28.100 168.200 28.200 ;
        RECT 187.800 28.100 188.200 28.200 ;
        RECT 192.600 28.100 193.000 28.200 ;
        RECT 167.800 27.800 193.000 28.100 ;
        RECT 13.400 26.800 13.800 27.200 ;
        RECT 25.400 27.100 25.800 27.200 ;
        RECT 35.800 27.100 36.100 27.800 ;
        RECT 61.400 27.200 61.700 27.800 ;
        RECT 25.400 26.800 36.100 27.100 ;
        RECT 39.800 27.100 40.200 27.200 ;
        RECT 45.400 27.100 45.800 27.200 ;
        RECT 47.800 27.100 48.200 27.200 ;
        RECT 39.800 26.800 48.200 27.100 ;
        RECT 55.800 26.800 56.200 27.200 ;
        RECT 61.400 26.800 61.800 27.200 ;
        RECT 63.000 27.100 63.400 27.200 ;
        RECT 65.400 27.100 65.800 27.200 ;
        RECT 69.400 27.100 69.800 27.200 ;
        RECT 63.000 26.800 69.800 27.100 ;
        RECT 71.800 26.800 72.200 27.200 ;
        RECT 76.600 26.800 77.000 27.200 ;
        RECT 79.800 27.100 80.200 27.200 ;
        RECT 83.000 27.100 83.300 27.800 ;
        RECT 95.000 27.200 95.300 27.800 ;
        RECT 104.600 27.200 104.900 27.800 ;
        RECT 111.800 27.200 112.100 27.800 ;
        RECT 84.600 27.100 85.000 27.200 ;
        RECT 79.800 26.800 85.000 27.100 ;
        RECT 86.200 27.100 86.600 27.200 ;
        RECT 90.200 27.100 90.600 27.200 ;
        RECT 86.200 26.800 90.600 27.100 ;
        RECT 91.000 27.100 91.400 27.200 ;
        RECT 91.800 27.100 92.200 27.200 ;
        RECT 91.000 26.800 92.200 27.100 ;
        RECT 92.600 27.100 93.000 27.200 ;
        RECT 94.200 27.100 94.600 27.200 ;
        RECT 92.600 26.800 94.600 27.100 ;
        RECT 95.000 26.800 95.400 27.200 ;
        RECT 95.800 27.100 96.200 27.200 ;
        RECT 96.600 27.100 97.000 27.200 ;
        RECT 95.800 26.800 97.000 27.100 ;
        RECT 97.400 26.800 97.800 27.200 ;
        RECT 98.200 26.800 98.600 27.200 ;
        RECT 104.600 26.800 105.000 27.200 ;
        RECT 109.400 27.100 109.800 27.200 ;
        RECT 111.800 27.100 112.200 27.200 ;
        RECT 109.400 26.800 112.200 27.100 ;
        RECT 113.400 27.100 113.800 27.200 ;
        RECT 116.600 27.100 117.000 27.200 ;
        RECT 113.400 26.800 117.000 27.100 ;
        RECT 117.400 27.100 117.700 27.800 ;
        RECT 125.400 27.100 125.800 27.200 ;
        RECT 117.400 26.800 125.800 27.100 ;
        RECT 127.800 27.100 128.200 27.200 ;
        RECT 133.400 27.100 133.800 27.200 ;
        RECT 146.200 27.100 146.600 27.200 ;
        RECT 127.800 26.800 133.800 27.100 ;
        RECT 140.600 26.800 146.600 27.100 ;
        RECT 147.800 27.100 148.200 27.200 ;
        RECT 155.800 27.100 156.200 27.200 ;
        RECT 160.600 27.100 161.000 27.200 ;
        RECT 179.800 27.100 180.200 27.200 ;
        RECT 147.800 26.800 180.200 27.100 ;
        RECT 180.600 26.800 181.000 27.200 ;
        RECT 181.400 27.100 181.800 27.200 ;
        RECT 190.200 27.100 190.600 27.200 ;
        RECT 198.200 27.100 198.600 27.200 ;
        RECT 181.400 26.800 198.600 27.100 ;
        RECT 6.200 26.100 6.600 26.200 ;
        RECT 13.400 26.100 13.700 26.800 ;
        RECT 55.800 26.200 56.100 26.800 ;
        RECT 6.200 25.800 13.700 26.100 ;
        RECT 22.200 26.100 22.600 26.200 ;
        RECT 32.600 26.100 33.000 26.200 ;
        RECT 46.200 26.100 46.600 26.200 ;
        RECT 22.200 25.800 46.600 26.100 ;
        RECT 54.200 26.100 54.600 26.200 ;
        RECT 55.000 26.100 55.400 26.200 ;
        RECT 54.200 25.800 55.400 26.100 ;
        RECT 55.800 25.800 56.200 26.200 ;
        RECT 59.000 26.100 59.400 26.200 ;
        RECT 71.800 26.100 72.100 26.800 ;
        RECT 76.600 26.200 76.900 26.800 ;
        RECT 59.000 25.800 72.100 26.100 ;
        RECT 72.600 26.100 73.000 26.200 ;
        RECT 73.400 26.100 73.800 26.200 ;
        RECT 72.600 25.800 73.800 26.100 ;
        RECT 76.600 25.800 77.000 26.200 ;
        RECT 83.000 26.100 83.400 26.200 ;
        RECT 88.600 26.100 89.000 26.200 ;
        RECT 89.400 26.100 89.800 26.200 ;
        RECT 83.000 25.800 88.100 26.100 ;
        RECT 88.600 25.800 89.800 26.100 ;
        RECT 93.400 26.100 93.800 26.200 ;
        RECT 97.400 26.100 97.700 26.800 ;
        RECT 93.400 25.800 97.700 26.100 ;
        RECT 98.200 26.200 98.500 26.800 ;
        RECT 140.600 26.200 140.900 26.800 ;
        RECT 98.200 25.800 98.600 26.200 ;
        RECT 99.800 26.100 100.200 26.200 ;
        RECT 100.600 26.100 101.000 26.200 ;
        RECT 99.800 25.800 101.000 26.100 ;
        RECT 103.800 26.100 104.200 26.200 ;
        RECT 113.400 26.100 113.800 26.200 ;
        RECT 103.800 25.800 113.800 26.100 ;
        RECT 114.200 26.100 114.600 26.200 ;
        RECT 120.600 26.100 121.000 26.200 ;
        RECT 114.200 25.800 121.000 26.100 ;
        RECT 123.800 26.100 124.200 26.200 ;
        RECT 124.600 26.100 125.000 26.200 ;
        RECT 123.800 25.800 125.000 26.100 ;
        RECT 127.000 26.100 127.400 26.200 ;
        RECT 131.800 26.100 132.200 26.200 ;
        RECT 127.000 25.800 132.200 26.100 ;
        RECT 140.600 25.800 141.000 26.200 ;
        RECT 144.600 26.100 145.000 26.200 ;
        RECT 156.600 26.100 157.000 26.200 ;
        RECT 144.600 25.800 157.000 26.100 ;
        RECT 163.800 26.100 164.200 26.200 ;
        RECT 164.600 26.100 165.000 26.200 ;
        RECT 163.800 25.800 165.000 26.100 ;
        RECT 175.800 26.100 176.200 26.200 ;
        RECT 180.600 26.100 180.900 26.800 ;
        RECT 175.800 25.800 180.900 26.100 ;
        RECT 192.600 26.100 193.000 26.200 ;
        RECT 199.800 26.100 200.200 26.200 ;
        RECT 203.000 26.100 203.400 26.200 ;
        RECT 192.600 25.800 203.400 26.100 ;
        RECT 87.800 25.200 88.100 25.800 ;
        RECT 38.200 25.100 38.600 25.200 ;
        RECT 48.600 25.100 49.000 25.200 ;
        RECT 50.200 25.100 50.600 25.200 ;
        RECT 38.200 24.800 45.700 25.100 ;
        RECT 48.600 24.800 50.600 25.100 ;
        RECT 61.400 25.100 61.800 25.200 ;
        RECT 63.000 25.100 63.400 25.200 ;
        RECT 72.600 25.100 73.000 25.200 ;
        RECT 74.200 25.100 74.600 25.200 ;
        RECT 61.400 24.800 63.400 25.100 ;
        RECT 65.400 24.800 70.500 25.100 ;
        RECT 71.800 24.800 74.600 25.100 ;
        RECT 87.800 24.800 88.200 25.200 ;
        RECT 90.200 25.100 90.600 25.200 ;
        RECT 112.600 25.100 113.000 25.200 ;
        RECT 118.200 25.100 118.600 25.200 ;
        RECT 90.200 24.800 118.600 25.100 ;
        RECT 120.600 25.100 121.000 25.200 ;
        RECT 122.200 25.100 122.600 25.200 ;
        RECT 124.600 25.100 125.000 25.200 ;
        RECT 120.600 24.800 125.000 25.100 ;
        RECT 162.200 25.100 162.600 25.200 ;
        RECT 163.800 25.100 164.200 25.200 ;
        RECT 162.200 24.800 164.200 25.100 ;
        RECT 167.800 25.100 168.200 25.200 ;
        RECT 186.200 25.100 186.600 25.200 ;
        RECT 194.200 25.100 194.600 25.200 ;
        RECT 167.800 24.800 194.600 25.100 ;
        RECT 45.400 24.200 45.700 24.800 ;
        RECT 65.400 24.200 65.700 24.800 ;
        RECT 70.200 24.200 70.500 24.800 ;
        RECT 45.400 23.800 45.800 24.200 ;
        RECT 65.400 23.800 65.800 24.200 ;
        RECT 70.200 23.800 70.600 24.200 ;
        RECT 77.400 24.100 77.800 24.200 ;
        RECT 103.800 24.100 104.200 24.200 ;
        RECT 77.400 23.800 104.200 24.100 ;
        RECT 126.200 24.100 126.600 24.200 ;
        RECT 130.200 24.100 130.600 24.200 ;
        RECT 126.200 23.800 130.600 24.100 ;
        RECT 15.000 23.100 15.400 23.200 ;
        RECT 59.800 23.100 60.200 23.200 ;
        RECT 15.000 22.800 60.200 23.100 ;
        RECT 60.600 23.100 61.000 23.200 ;
        RECT 62.200 23.100 62.600 23.200 ;
        RECT 60.600 22.800 62.600 23.100 ;
        RECT 68.600 23.100 69.000 23.200 ;
        RECT 81.400 23.100 81.800 23.200 ;
        RECT 68.600 22.800 81.800 23.100 ;
        RECT 104.600 23.100 105.000 23.200 ;
        RECT 106.200 23.100 106.600 23.200 ;
        RECT 104.600 22.800 106.600 23.100 ;
        RECT 118.200 22.800 118.600 23.200 ;
        RECT 119.000 23.100 119.400 23.200 ;
        RECT 182.200 23.100 182.600 23.200 ;
        RECT 119.000 22.800 182.600 23.100 ;
        RECT 62.200 22.100 62.600 22.200 ;
        RECT 66.200 22.100 66.600 22.200 ;
        RECT 78.200 22.100 78.600 22.200 ;
        RECT 62.200 21.800 78.600 22.100 ;
        RECT 79.800 21.800 80.200 22.200 ;
        RECT 87.000 22.100 87.400 22.200 ;
        RECT 94.200 22.100 94.600 22.200 ;
        RECT 118.200 22.100 118.500 22.800 ;
        RECT 87.000 21.800 89.700 22.100 ;
        RECT 94.200 21.800 118.500 22.100 ;
        RECT 195.800 22.100 196.200 22.200 ;
        RECT 199.000 22.100 199.400 22.200 ;
        RECT 195.800 21.800 199.400 22.100 ;
        RECT 79.800 21.200 80.100 21.800 ;
        RECT 89.400 21.200 89.700 21.800 ;
        RECT 79.800 20.800 80.200 21.200 ;
        RECT 89.400 20.800 89.800 21.200 ;
        RECT 94.200 21.100 94.600 21.200 ;
        RECT 100.600 21.100 101.000 21.200 ;
        RECT 94.200 20.800 101.000 21.100 ;
        RECT 115.800 21.100 116.200 21.200 ;
        RECT 127.800 21.100 128.200 21.200 ;
        RECT 129.400 21.100 129.800 21.200 ;
        RECT 115.800 20.800 129.800 21.100 ;
        RECT 81.400 20.100 81.800 20.200 ;
        RECT 114.200 20.100 114.600 20.200 ;
        RECT 81.400 19.800 114.600 20.100 ;
        RECT 38.200 19.100 38.600 19.200 ;
        RECT 67.800 19.100 68.200 19.200 ;
        RECT 37.400 18.800 68.200 19.100 ;
        RECT 69.400 19.100 69.800 19.200 ;
        RECT 88.600 19.100 89.000 19.200 ;
        RECT 69.400 18.800 89.000 19.100 ;
        RECT 95.800 19.100 96.200 19.200 ;
        RECT 163.800 19.100 164.200 19.200 ;
        RECT 95.800 18.800 164.200 19.100 ;
        RECT 195.000 19.100 195.400 19.200 ;
        RECT 195.000 18.800 196.900 19.100 ;
        RECT 196.600 18.200 196.900 18.800 ;
        RECT 31.800 17.800 32.200 18.200 ;
        RECT 50.200 18.100 50.600 18.200 ;
        RECT 56.600 18.100 57.000 18.200 ;
        RECT 50.200 17.800 57.000 18.100 ;
        RECT 102.200 18.100 102.600 18.200 ;
        RECT 142.200 18.100 142.600 18.200 ;
        RECT 146.200 18.100 146.600 18.200 ;
        RECT 102.200 17.800 146.600 18.100 ;
        RECT 159.800 18.100 160.200 18.200 ;
        RECT 160.600 18.100 161.000 18.200 ;
        RECT 162.200 18.100 162.600 18.200 ;
        RECT 178.200 18.100 178.600 18.200 ;
        RECT 180.600 18.100 181.000 18.200 ;
        RECT 159.800 17.800 181.000 18.100 ;
        RECT 196.600 17.800 197.000 18.200 ;
        RECT 31.800 17.200 32.100 17.800 ;
        RECT 25.400 17.100 25.800 17.200 ;
        RECT 30.200 17.100 30.600 17.200 ;
        RECT 25.400 16.800 30.600 17.100 ;
        RECT 31.800 16.800 32.200 17.200 ;
        RECT 34.200 17.100 34.600 17.200 ;
        RECT 51.800 17.100 52.200 17.200 ;
        RECT 55.000 17.100 55.400 17.200 ;
        RECT 34.200 16.800 55.400 17.100 ;
        RECT 65.400 17.100 65.800 17.200 ;
        RECT 67.800 17.100 68.200 17.200 ;
        RECT 72.600 17.100 73.000 17.200 ;
        RECT 65.400 16.800 73.000 17.100 ;
        RECT 87.800 16.800 88.200 17.200 ;
        RECT 88.600 17.100 89.000 17.200 ;
        RECT 100.600 17.100 101.000 17.200 ;
        RECT 111.000 17.100 111.400 17.200 ;
        RECT 88.600 16.800 111.400 17.100 ;
        RECT 115.000 17.100 115.400 17.200 ;
        RECT 115.800 17.100 116.200 17.200 ;
        RECT 115.000 16.800 116.200 17.100 ;
        RECT 141.400 17.100 141.800 17.200 ;
        RECT 146.200 17.100 146.600 17.200 ;
        RECT 155.800 17.100 156.200 17.200 ;
        RECT 141.400 16.800 156.200 17.100 ;
        RECT 163.000 17.100 163.400 17.200 ;
        RECT 168.600 17.100 169.000 17.200 ;
        RECT 185.400 17.100 185.800 17.200 ;
        RECT 187.000 17.100 187.400 17.200 ;
        RECT 163.000 16.800 187.400 17.100 ;
        RECT 87.800 16.200 88.100 16.800 ;
        RECT 10.200 16.100 10.600 16.200 ;
        RECT 11.800 16.100 12.200 16.200 ;
        RECT 10.200 15.800 12.200 16.100 ;
        RECT 26.200 16.100 26.600 16.200 ;
        RECT 29.400 16.100 29.800 16.200 ;
        RECT 86.200 16.100 86.600 16.200 ;
        RECT 87.800 16.100 88.200 16.200 ;
        RECT 26.200 15.800 88.200 16.100 ;
        RECT 107.000 16.100 107.400 16.200 ;
        RECT 115.000 16.100 115.400 16.200 ;
        RECT 107.000 15.800 115.400 16.100 ;
        RECT 117.400 16.100 117.800 16.200 ;
        RECT 122.200 16.100 122.600 16.200 ;
        RECT 117.400 15.800 122.600 16.100 ;
        RECT 136.600 16.100 137.000 16.200 ;
        RECT 165.400 16.100 165.800 16.200 ;
        RECT 136.600 15.800 165.800 16.100 ;
        RECT 11.000 15.100 11.400 15.200 ;
        RECT 14.200 15.100 14.600 15.200 ;
        RECT 18.200 15.100 18.600 15.200 ;
        RECT 11.000 14.800 18.600 15.100 ;
        RECT 19.800 15.100 20.200 15.200 ;
        RECT 27.800 15.100 28.200 15.200 ;
        RECT 19.800 14.800 28.200 15.100 ;
        RECT 31.800 15.100 32.200 15.200 ;
        RECT 34.200 15.100 34.600 15.200 ;
        RECT 31.800 14.800 34.600 15.100 ;
        RECT 44.600 15.100 45.000 15.200 ;
        RECT 61.400 15.100 61.800 15.200 ;
        RECT 79.800 15.100 80.200 15.200 ;
        RECT 99.800 15.100 100.200 15.200 ;
        RECT 44.600 14.800 53.700 15.100 ;
        RECT 61.400 14.800 79.300 15.100 ;
        RECT 79.800 14.800 100.200 15.100 ;
        RECT 115.800 15.100 116.200 15.200 ;
        RECT 119.000 15.100 119.400 15.200 ;
        RECT 115.800 14.800 119.400 15.100 ;
        RECT 173.400 15.100 173.800 15.200 ;
        RECT 183.000 15.100 183.400 15.200 ;
        RECT 186.200 15.100 186.600 15.200 ;
        RECT 173.400 14.800 186.600 15.100 ;
        RECT 53.400 14.200 53.700 14.800 ;
        RECT 9.400 14.100 9.800 14.200 ;
        RECT 15.000 14.100 15.400 14.200 ;
        RECT 9.400 13.800 15.400 14.100 ;
        RECT 26.200 14.100 26.600 14.200 ;
        RECT 31.800 14.100 32.200 14.200 ;
        RECT 32.600 14.100 33.000 14.200 ;
        RECT 26.200 13.800 33.000 14.100 ;
        RECT 36.600 14.100 37.000 14.200 ;
        RECT 38.200 14.100 38.600 14.200 ;
        RECT 43.000 14.100 43.400 14.200 ;
        RECT 36.600 13.800 43.400 14.100 ;
        RECT 53.400 13.800 53.800 14.200 ;
        RECT 71.800 14.100 72.200 14.200 ;
        RECT 72.600 14.100 73.000 14.200 ;
        RECT 71.800 13.800 73.000 14.100 ;
        RECT 79.000 14.100 79.300 14.800 ;
        RECT 82.200 14.100 82.600 14.200 ;
        RECT 79.000 13.800 82.600 14.100 ;
        RECT 98.200 13.800 98.600 14.200 ;
        RECT 118.200 14.100 118.600 14.200 ;
        RECT 119.000 14.100 119.400 14.200 ;
        RECT 118.200 13.800 119.400 14.100 ;
        RECT 125.400 13.800 125.800 14.200 ;
        RECT 143.000 14.100 143.400 14.200 ;
        RECT 146.200 14.100 146.600 14.200 ;
        RECT 159.800 14.100 160.200 14.200 ;
        RECT 143.000 13.800 160.200 14.100 ;
        RECT 163.000 13.800 163.400 14.200 ;
        RECT 165.400 14.100 165.800 14.200 ;
        RECT 167.800 14.100 168.200 14.200 ;
        RECT 165.400 13.800 168.200 14.100 ;
        RECT 5.400 13.100 5.800 13.200 ;
        RECT 11.000 13.100 11.400 13.200 ;
        RECT 5.400 12.800 11.400 13.100 ;
        RECT 35.800 13.100 36.200 13.200 ;
        RECT 39.000 13.100 39.400 13.200 ;
        RECT 35.800 12.800 39.400 13.100 ;
        RECT 39.800 13.100 40.200 13.200 ;
        RECT 41.400 13.100 41.800 13.200 ;
        RECT 39.800 12.800 41.800 13.100 ;
        RECT 74.200 13.100 74.600 13.200 ;
        RECT 79.000 13.100 79.400 13.200 ;
        RECT 74.200 12.800 79.400 13.100 ;
        RECT 98.200 13.100 98.500 13.800 ;
        RECT 99.000 13.100 99.400 13.200 ;
        RECT 98.200 12.800 99.400 13.100 ;
        RECT 110.200 13.100 110.600 13.200 ;
        RECT 114.200 13.100 114.600 13.200 ;
        RECT 125.400 13.100 125.700 13.800 ;
        RECT 163.000 13.200 163.300 13.800 ;
        RECT 151.000 13.100 151.400 13.200 ;
        RECT 110.200 12.800 125.700 13.100 ;
        RECT 144.600 12.800 151.400 13.100 ;
        RECT 163.000 12.800 163.400 13.200 ;
        RECT 144.600 12.200 144.900 12.800 ;
        RECT 26.200 11.800 26.600 12.200 ;
        RECT 39.000 12.100 39.400 12.200 ;
        RECT 57.400 12.100 57.800 12.200 ;
        RECT 39.000 11.800 57.800 12.100 ;
        RECT 110.200 12.100 110.600 12.200 ;
        RECT 120.600 12.100 121.000 12.200 ;
        RECT 110.200 11.800 121.000 12.100 ;
        RECT 144.600 11.800 145.000 12.200 ;
        RECT 186.200 12.100 186.600 12.200 ;
        RECT 187.000 12.100 187.400 12.200 ;
        RECT 186.200 11.800 187.400 12.100 ;
        RECT 26.200 11.200 26.500 11.800 ;
        RECT 26.200 11.100 26.600 11.200 ;
        RECT 28.600 11.100 29.000 11.200 ;
        RECT 26.200 10.800 29.000 11.100 ;
        RECT 68.600 11.100 69.000 11.200 ;
        RECT 84.600 11.100 85.000 11.200 ;
        RECT 68.600 10.800 85.000 11.100 ;
        RECT 163.800 11.100 164.200 11.200 ;
        RECT 173.400 11.100 173.800 11.200 ;
        RECT 176.600 11.100 177.000 11.200 ;
        RECT 163.800 10.800 177.000 11.100 ;
        RECT 24.600 10.100 25.000 10.200 ;
        RECT 75.800 10.100 76.200 10.200 ;
        RECT 24.600 9.800 76.200 10.100 ;
        RECT 83.800 10.100 84.200 10.200 ;
        RECT 86.200 10.100 86.600 10.200 ;
        RECT 91.000 10.100 91.400 10.200 ;
        RECT 83.800 9.800 91.400 10.100 ;
        RECT 157.400 10.100 157.800 10.200 ;
        RECT 162.200 10.100 162.600 10.200 ;
        RECT 157.400 9.800 162.600 10.100 ;
        RECT 28.600 9.100 29.000 9.200 ;
        RECT 41.400 9.100 41.800 9.200 ;
        RECT 87.800 9.100 88.200 9.200 ;
        RECT 28.600 8.800 88.200 9.100 ;
        RECT 103.000 9.100 103.400 9.200 ;
        RECT 103.800 9.100 104.200 9.200 ;
        RECT 111.800 9.100 112.200 9.200 ;
        RECT 103.000 8.800 112.200 9.100 ;
        RECT 115.000 9.100 115.400 9.200 ;
        RECT 119.000 9.100 119.400 9.200 ;
        RECT 122.200 9.100 122.600 9.200 ;
        RECT 115.000 8.800 122.600 9.100 ;
        RECT 131.000 9.100 131.400 9.200 ;
        RECT 133.400 9.100 133.800 9.200 ;
        RECT 137.400 9.100 137.800 9.200 ;
        RECT 131.000 8.800 137.800 9.100 ;
        RECT 153.400 9.100 153.800 9.200 ;
        RECT 156.600 9.100 157.000 9.200 ;
        RECT 153.400 8.800 157.000 9.100 ;
        RECT 159.000 9.100 159.400 9.200 ;
        RECT 161.400 9.100 161.800 9.200 ;
        RECT 159.000 8.800 161.800 9.100 ;
        RECT 198.200 9.100 198.600 9.200 ;
        RECT 202.200 9.100 202.600 9.200 ;
        RECT 198.200 8.800 202.600 9.100 ;
        RECT 29.400 8.100 29.800 8.200 ;
        RECT 68.600 8.100 69.000 8.200 ;
        RECT 29.400 7.800 69.000 8.100 ;
        RECT 70.200 7.800 70.600 8.200 ;
        RECT 78.200 8.100 78.600 8.200 ;
        RECT 80.600 8.100 81.000 8.200 ;
        RECT 78.200 7.800 81.000 8.100 ;
        RECT 107.800 8.100 108.200 8.200 ;
        RECT 116.600 8.100 117.000 8.200 ;
        RECT 107.800 7.800 117.000 8.100 ;
        RECT 121.400 7.800 121.800 8.200 ;
        RECT 131.000 7.800 131.400 8.200 ;
        RECT 160.600 7.800 161.000 8.200 ;
        RECT 171.800 7.800 172.200 8.200 ;
        RECT 59.800 7.100 60.200 7.200 ;
        RECT 70.200 7.100 70.500 7.800 ;
        RECT 121.400 7.200 121.700 7.800 ;
        RECT 84.600 7.100 85.000 7.200 ;
        RECT 91.800 7.100 92.200 7.200 ;
        RECT 94.200 7.100 94.600 7.200 ;
        RECT 105.400 7.100 105.800 7.200 ;
        RECT 14.200 6.800 31.300 7.100 ;
        RECT 59.800 6.800 105.800 7.100 ;
        RECT 108.600 6.800 109.000 7.200 ;
        RECT 117.400 7.100 117.800 7.200 ;
        RECT 121.400 7.100 121.800 7.200 ;
        RECT 117.400 6.800 121.800 7.100 ;
        RECT 131.000 7.100 131.300 7.800 ;
        RECT 137.400 7.100 137.800 7.200 ;
        RECT 131.000 6.800 137.800 7.100 ;
        RECT 160.600 7.100 160.900 7.800 ;
        RECT 171.800 7.100 172.100 7.800 ;
        RECT 176.600 7.100 177.000 7.200 ;
        RECT 186.200 7.100 186.600 7.200 ;
        RECT 160.600 6.800 186.600 7.100 ;
        RECT 14.200 6.200 14.500 6.800 ;
        RECT 15.800 6.200 16.100 6.800 ;
        RECT 31.000 6.200 31.300 6.800 ;
        RECT 14.200 5.800 14.600 6.200 ;
        RECT 15.800 5.800 16.200 6.200 ;
        RECT 19.000 6.100 19.400 6.200 ;
        RECT 27.000 6.100 27.400 6.200 ;
        RECT 19.000 5.800 27.400 6.100 ;
        RECT 28.600 6.100 29.000 6.200 ;
        RECT 29.400 6.100 29.800 6.200 ;
        RECT 28.600 5.800 29.800 6.100 ;
        RECT 31.000 6.100 31.400 6.200 ;
        RECT 43.800 6.100 44.200 6.200 ;
        RECT 47.000 6.100 47.400 6.200 ;
        RECT 31.000 5.800 47.400 6.100 ;
        RECT 58.200 6.100 58.600 6.200 ;
        RECT 65.400 6.100 65.800 6.200 ;
        RECT 58.200 5.800 65.800 6.100 ;
        RECT 86.200 6.100 86.600 6.200 ;
        RECT 95.800 6.100 96.200 6.200 ;
        RECT 86.200 5.800 96.200 6.100 ;
        RECT 108.600 6.100 108.900 6.800 ;
        RECT 113.400 6.100 113.800 6.200 ;
        RECT 108.600 5.800 113.800 6.100 ;
        RECT 116.600 6.100 117.000 6.200 ;
        RECT 121.400 6.100 121.800 6.200 ;
        RECT 116.600 5.800 121.800 6.100 ;
        RECT 48.600 5.100 49.000 5.200 ;
        RECT 41.400 4.800 49.000 5.100 ;
        RECT 66.200 5.100 66.600 5.200 ;
        RECT 67.800 5.100 68.200 5.200 ;
        RECT 78.200 5.100 78.600 5.200 ;
        RECT 112.600 5.100 113.000 5.200 ;
        RECT 115.800 5.100 116.200 5.200 ;
        RECT 66.200 4.800 116.200 5.100 ;
        RECT 120.600 5.100 121.000 5.200 ;
        RECT 127.000 5.100 127.400 5.200 ;
        RECT 120.600 4.800 127.400 5.100 ;
        RECT 41.400 4.200 41.700 4.800 ;
        RECT 41.400 3.800 41.800 4.200 ;
      LAYER via3 ;
        RECT 196.600 176.800 197.000 177.200 ;
        RECT 111.800 171.800 112.200 172.200 ;
        RECT 48.600 169.800 49.000 170.200 ;
        RECT 106.200 167.800 106.600 168.200 ;
        RECT 155.000 166.800 155.400 167.200 ;
        RECT 190.200 166.800 190.600 167.200 ;
        RECT 112.600 165.800 113.000 166.200 ;
        RECT 66.200 164.800 66.600 165.200 ;
        RECT 71.800 163.800 72.200 164.200 ;
        RECT 197.400 163.800 197.800 164.200 ;
        RECT 73.400 162.800 73.800 163.200 ;
        RECT 77.400 159.800 77.800 160.200 ;
        RECT 84.600 158.800 85.000 159.200 ;
        RECT 21.400 155.800 21.800 156.200 ;
        RECT 151.800 153.800 152.200 154.200 ;
        RECT 190.200 153.800 190.600 154.200 ;
        RECT 14.200 152.800 14.600 153.200 ;
        RECT 138.200 152.800 138.600 153.200 ;
        RECT 175.000 152.800 175.400 153.200 ;
        RECT 61.400 150.800 61.800 151.200 ;
        RECT 196.600 150.800 197.000 151.200 ;
        RECT 39.000 149.800 39.400 150.200 ;
        RECT 125.400 149.800 125.800 150.200 ;
        RECT 62.200 148.800 62.600 149.200 ;
        RECT 25.400 147.800 25.800 148.200 ;
        RECT 84.600 147.800 85.000 148.200 ;
        RECT 123.800 146.800 124.200 147.200 ;
        RECT 174.200 146.800 174.600 147.200 ;
        RECT 24.600 145.800 25.000 146.200 ;
        RECT 54.200 145.800 54.600 146.200 ;
        RECT 155.000 145.800 155.400 146.200 ;
        RECT 185.400 145.800 185.800 146.200 ;
        RECT 105.400 144.800 105.800 145.200 ;
        RECT 183.000 144.800 183.400 145.200 ;
        RECT 190.200 144.800 190.600 145.200 ;
        RECT 13.400 143.800 13.800 144.200 ;
        RECT 100.600 142.800 101.000 143.200 ;
        RECT 123.000 142.800 123.400 143.200 ;
        RECT 199.800 142.800 200.200 143.200 ;
        RECT 161.400 141.800 161.800 142.200 ;
        RECT 195.800 141.800 196.200 142.200 ;
        RECT 128.600 140.800 129.000 141.200 ;
        RECT 147.000 140.800 147.400 141.200 ;
        RECT 173.400 140.800 173.800 141.200 ;
        RECT 199.800 140.800 200.200 141.200 ;
        RECT 173.400 139.800 173.800 140.200 ;
        RECT 21.400 138.800 21.800 139.200 ;
        RECT 127.800 138.800 128.200 139.200 ;
        RECT 127.000 136.800 127.400 137.200 ;
        RECT 164.600 136.800 165.000 137.200 ;
        RECT 120.600 135.800 121.000 136.200 ;
        RECT 199.000 135.800 199.400 136.200 ;
        RECT 19.000 134.800 19.400 135.200 ;
        RECT 123.000 134.800 123.400 135.200 ;
        RECT 128.600 133.800 129.000 134.200 ;
        RECT 179.000 133.800 179.400 134.200 ;
        RECT 80.600 132.800 81.000 133.200 ;
        RECT 165.400 132.800 165.800 133.200 ;
        RECT 82.200 131.800 82.600 132.200 ;
        RECT 135.800 131.800 136.200 132.200 ;
        RECT 41.400 130.800 41.800 131.200 ;
        RECT 43.800 130.800 44.200 131.200 ;
        RECT 115.000 130.800 115.400 131.200 ;
        RECT 196.600 129.800 197.000 130.200 ;
        RECT 89.400 128.800 89.800 129.200 ;
        RECT 40.600 127.800 41.000 128.200 ;
        RECT 103.800 126.800 104.200 127.200 ;
        RECT 139.000 126.800 139.400 127.200 ;
        RECT 34.200 125.800 34.600 126.200 ;
        RECT 139.800 125.800 140.200 126.200 ;
        RECT 183.800 124.800 184.200 125.200 ;
        RECT 113.400 123.800 113.800 124.200 ;
        RECT 171.000 123.800 171.400 124.200 ;
        RECT 53.400 122.800 53.800 123.200 ;
        RECT 76.600 121.800 77.000 122.200 ;
        RECT 81.400 120.800 81.800 121.200 ;
        RECT 173.400 120.800 173.800 121.200 ;
        RECT 64.600 117.800 65.000 118.200 ;
        RECT 86.200 117.800 86.600 118.200 ;
        RECT 58.200 116.800 58.600 117.200 ;
        RECT 65.400 115.800 65.800 116.200 ;
        RECT 92.600 115.800 93.000 116.200 ;
        RECT 145.400 115.800 145.800 116.200 ;
        RECT 157.400 115.800 157.800 116.200 ;
        RECT 42.200 114.800 42.600 115.200 ;
        RECT 99.800 114.800 100.200 115.200 ;
        RECT 160.600 114.800 161.000 115.200 ;
        RECT 54.200 113.800 54.600 114.200 ;
        RECT 67.800 112.800 68.200 113.200 ;
        RECT 146.200 112.800 146.600 113.200 ;
        RECT 194.200 111.800 194.600 112.200 ;
        RECT 48.600 110.800 49.000 111.200 ;
        RECT 151.000 109.800 151.400 110.200 ;
        RECT 193.400 109.800 193.800 110.200 ;
        RECT 72.600 107.800 73.000 108.200 ;
        RECT 170.200 107.800 170.600 108.200 ;
        RECT 17.400 106.800 17.800 107.200 ;
        RECT 54.200 106.800 54.600 107.200 ;
        RECT 41.400 105.800 41.800 106.200 ;
        RECT 192.600 105.800 193.000 106.200 ;
        RECT 69.400 104.800 69.800 105.200 ;
        RECT 43.800 103.800 44.200 104.200 ;
        RECT 121.400 103.800 121.800 104.200 ;
        RECT 89.400 100.800 89.800 101.200 ;
        RECT 191.000 100.800 191.400 101.200 ;
        RECT 76.600 99.800 77.000 100.200 ;
        RECT 92.600 97.800 93.000 98.200 ;
        RECT 53.400 96.800 53.800 97.200 ;
        RECT 72.600 96.800 73.000 97.200 ;
        RECT 22.200 95.800 22.600 96.200 ;
        RECT 39.800 95.800 40.200 96.200 ;
        RECT 64.600 94.800 65.000 95.200 ;
        RECT 83.000 94.800 83.400 95.200 ;
        RECT 139.000 94.800 139.400 95.200 ;
        RECT 46.200 93.800 46.600 94.200 ;
        RECT 59.800 93.800 60.200 94.200 ;
        RECT 79.800 93.800 80.200 94.200 ;
        RECT 162.200 93.800 162.600 94.200 ;
        RECT 40.600 92.800 41.000 93.200 ;
        RECT 85.400 92.800 85.800 93.200 ;
        RECT 90.200 92.800 90.600 93.200 ;
        RECT 31.000 91.800 31.400 92.200 ;
        RECT 80.600 91.800 81.000 92.200 ;
        RECT 115.800 91.800 116.200 92.200 ;
        RECT 37.400 90.800 37.800 91.200 ;
        RECT 75.800 90.800 76.200 91.200 ;
        RECT 159.800 90.800 160.200 91.200 ;
        RECT 32.600 88.800 33.000 89.200 ;
        RECT 65.400 88.800 65.800 89.200 ;
        RECT 70.200 88.800 70.600 89.200 ;
        RECT 83.800 88.800 84.200 89.200 ;
        RECT 147.800 88.800 148.200 89.200 ;
        RECT 65.400 87.800 65.800 88.200 ;
        RECT 44.600 86.800 45.000 87.200 ;
        RECT 99.000 86.800 99.400 87.200 ;
        RECT 13.400 85.800 13.800 86.200 ;
        RECT 75.000 85.800 75.400 86.200 ;
        RECT 78.200 85.800 78.600 86.200 ;
        RECT 82.200 85.800 82.600 86.200 ;
        RECT 87.000 85.800 87.400 86.200 ;
        RECT 195.000 85.800 195.400 86.200 ;
        RECT 201.400 85.800 201.800 86.200 ;
        RECT 162.200 84.800 162.600 85.200 ;
        RECT 60.600 83.800 61.000 84.200 ;
        RECT 159.000 83.800 159.400 84.200 ;
        RECT 58.200 82.800 58.600 83.200 ;
        RECT 168.600 82.800 169.000 83.200 ;
        RECT 95.000 81.800 95.400 82.200 ;
        RECT 13.400 80.800 13.800 81.200 ;
        RECT 18.200 80.800 18.600 81.200 ;
        RECT 47.000 80.800 47.400 81.200 ;
        RECT 77.400 78.800 77.800 79.200 ;
        RECT 119.000 78.800 119.400 79.200 ;
        RECT 100.600 77.800 101.000 78.200 ;
        RECT 52.600 76.800 53.000 77.200 ;
        RECT 99.000 76.800 99.400 77.200 ;
        RECT 140.600 76.800 141.000 77.200 ;
        RECT 47.000 75.800 47.400 76.200 ;
        RECT 49.400 75.800 49.800 76.200 ;
        RECT 107.000 75.800 107.400 76.200 ;
        RECT 115.000 75.800 115.400 76.200 ;
        RECT 161.400 75.800 161.800 76.200 ;
        RECT 55.000 74.800 55.400 75.200 ;
        RECT 14.200 73.800 14.600 74.200 ;
        RECT 18.200 73.800 18.600 74.200 ;
        RECT 76.600 74.800 77.000 75.200 ;
        RECT 84.600 74.800 85.000 75.200 ;
        RECT 105.400 74.800 105.800 75.200 ;
        RECT 129.400 74.800 129.800 75.200 ;
        RECT 159.800 74.800 160.200 75.200 ;
        RECT 73.400 73.800 73.800 74.200 ;
        RECT 83.000 73.800 83.400 74.200 ;
        RECT 91.800 73.800 92.200 74.200 ;
        RECT 123.800 73.800 124.200 74.200 ;
        RECT 170.200 73.800 170.600 74.200 ;
        RECT 71.800 72.800 72.200 73.200 ;
        RECT 142.200 72.800 142.600 73.200 ;
        RECT 169.400 72.800 169.800 73.200 ;
        RECT 193.400 72.800 193.800 73.200 ;
        RECT 69.400 71.800 69.800 72.200 ;
        RECT 116.600 71.800 117.000 72.200 ;
        RECT 122.200 71.800 122.600 72.200 ;
        RECT 180.600 71.800 181.000 72.200 ;
        RECT 28.600 70.800 29.000 71.200 ;
        RECT 56.600 69.800 57.000 70.200 ;
        RECT 151.000 69.800 151.400 70.200 ;
        RECT 135.000 67.800 135.400 68.200 ;
        RECT 147.000 67.800 147.400 68.200 ;
        RECT 85.400 66.800 85.800 67.200 ;
        RECT 99.800 66.800 100.200 67.200 ;
        RECT 128.600 66.800 129.000 67.200 ;
        RECT 149.400 66.800 149.800 67.200 ;
        RECT 152.600 66.800 153.000 67.200 ;
        RECT 14.200 65.800 14.600 66.200 ;
        RECT 161.400 65.800 161.800 66.200 ;
        RECT 168.600 65.800 169.000 66.200 ;
        RECT 88.600 63.800 89.000 64.200 ;
        RECT 83.800 61.800 84.200 62.200 ;
        RECT 90.200 61.800 90.600 62.200 ;
        RECT 126.200 61.800 126.600 62.200 ;
        RECT 139.000 60.800 139.400 61.200 ;
        RECT 26.200 58.800 26.600 59.200 ;
        RECT 68.600 58.800 69.000 59.200 ;
        RECT 118.200 58.800 118.600 59.200 ;
        RECT 148.600 58.800 149.000 59.200 ;
        RECT 79.000 57.800 79.400 58.200 ;
        RECT 35.000 56.800 35.400 57.200 ;
        RECT 110.200 56.800 110.600 57.200 ;
        RECT 58.200 55.800 58.600 56.200 ;
        RECT 87.800 55.800 88.200 56.200 ;
        RECT 59.000 54.800 59.400 55.200 ;
        RECT 119.000 54.800 119.400 55.200 ;
        RECT 59.800 53.800 60.200 54.200 ;
        RECT 111.800 53.800 112.200 54.200 ;
        RECT 67.800 52.800 68.200 53.200 ;
        RECT 99.800 52.800 100.200 53.200 ;
        RECT 163.800 52.800 164.200 53.200 ;
        RECT 104.600 51.800 105.000 52.200 ;
        RECT 117.400 51.800 117.800 52.200 ;
        RECT 91.800 48.800 92.200 49.200 ;
        RECT 31.800 47.800 32.200 48.200 ;
        RECT 201.400 47.800 201.800 48.200 ;
        RECT 103.800 46.800 104.200 47.200 ;
        RECT 105.400 46.800 105.800 47.200 ;
        RECT 147.800 46.800 148.200 47.200 ;
        RECT 155.000 46.800 155.400 47.200 ;
        RECT 12.600 45.800 13.000 46.200 ;
        RECT 96.600 45.800 97.000 46.200 ;
        RECT 98.200 45.800 98.600 46.200 ;
        RECT 116.600 45.800 117.000 46.200 ;
        RECT 49.400 44.800 49.800 45.200 ;
        RECT 115.800 44.800 116.200 45.200 ;
        RECT 127.000 44.800 127.400 45.200 ;
        RECT 149.400 44.800 149.800 45.200 ;
        RECT 164.600 44.800 165.000 45.200 ;
        RECT 108.600 43.800 109.000 44.200 ;
        RECT 43.800 41.800 44.200 42.200 ;
        RECT 63.000 41.800 63.400 42.200 ;
        RECT 165.400 41.800 165.800 42.200 ;
        RECT 171.000 41.800 171.400 42.200 ;
        RECT 187.000 41.800 187.400 42.200 ;
        RECT 119.000 40.800 119.400 41.200 ;
        RECT 62.200 39.800 62.600 40.200 ;
        RECT 106.200 39.800 106.600 40.200 ;
        RECT 28.600 36.800 29.000 37.200 ;
        RECT 98.200 36.800 98.600 37.200 ;
        RECT 16.600 35.800 17.000 36.200 ;
        RECT 37.400 35.800 37.800 36.200 ;
        RECT 17.400 34.800 17.800 35.200 ;
        RECT 70.200 34.800 70.600 35.200 ;
        RECT 95.000 34.800 95.400 35.200 ;
        RECT 29.400 33.800 29.800 34.200 ;
        RECT 49.400 33.800 49.800 34.200 ;
        RECT 106.200 33.800 106.600 34.200 ;
        RECT 71.000 32.800 71.400 33.200 ;
        RECT 77.400 31.800 77.800 32.200 ;
        RECT 96.600 30.800 97.000 31.200 ;
        RECT 50.200 29.800 50.600 30.200 ;
        RECT 35.000 28.800 35.400 29.200 ;
        RECT 171.000 28.800 171.400 29.200 ;
        RECT 81.400 27.800 81.800 28.200 ;
        RECT 93.400 27.800 93.800 28.200 ;
        RECT 90.200 26.800 90.600 27.200 ;
        RECT 91.800 26.800 92.200 27.200 ;
        RECT 111.800 26.800 112.200 27.200 ;
        RECT 179.800 26.800 180.200 27.200 ;
        RECT 199.800 25.800 200.200 26.200 ;
        RECT 118.200 24.800 118.600 25.200 ;
        RECT 122.200 24.800 122.600 25.200 ;
        RECT 186.200 24.800 186.600 25.200 ;
        RECT 103.800 23.800 104.200 24.200 ;
        RECT 127.800 20.800 128.200 21.200 ;
        RECT 114.200 19.800 114.600 20.200 ;
        RECT 88.600 18.800 89.000 19.200 ;
        RECT 160.600 17.800 161.000 18.200 ;
        RECT 111.000 16.800 111.400 17.200 ;
        RECT 115.800 16.800 116.200 17.200 ;
        RECT 18.200 14.800 18.600 15.200 ;
        RECT 119.000 13.800 119.400 14.200 ;
        RECT 84.600 10.800 85.000 11.200 ;
        RECT 86.200 9.800 86.600 10.200 ;
        RECT 121.400 6.800 121.800 7.200 ;
        RECT 29.400 5.800 29.800 6.200 ;
      LAYER metal4 ;
        RECT 196.600 176.800 197.000 177.200 ;
        RECT 196.600 173.200 196.900 176.800 ;
        RECT 196.600 172.800 197.000 173.200 ;
        RECT 111.800 171.800 112.200 172.200 ;
        RECT 190.200 171.800 190.600 172.200 ;
        RECT 48.600 169.800 49.000 170.200 ;
        RECT 24.600 161.800 25.000 162.200 ;
        RECT 21.400 155.800 21.800 156.200 ;
        RECT 14.200 152.800 14.600 153.200 ;
        RECT 12.600 144.800 13.000 145.200 ;
        RECT 12.600 126.200 12.900 144.800 ;
        RECT 13.400 143.800 13.800 144.200 ;
        RECT 13.400 136.200 13.700 143.800 ;
        RECT 13.400 135.800 13.800 136.200 ;
        RECT 12.600 125.800 13.000 126.200 ;
        RECT 13.400 86.200 13.700 135.800 ;
        RECT 12.600 85.800 13.000 86.200 ;
        RECT 13.400 85.800 13.800 86.200 ;
        RECT 12.600 51.200 12.900 85.800 ;
        RECT 13.400 80.800 13.800 81.200 ;
        RECT 13.400 66.100 13.700 80.800 ;
        RECT 14.200 74.200 14.500 152.800 ;
        RECT 19.000 143.800 19.400 144.200 ;
        RECT 19.000 135.200 19.300 143.800 ;
        RECT 21.400 139.200 21.700 155.800 ;
        RECT 24.600 146.200 24.900 161.800 ;
        RECT 44.600 153.800 45.000 154.200 ;
        RECT 39.000 149.800 39.400 150.200 ;
        RECT 25.400 147.800 25.800 148.200 ;
        RECT 24.600 145.800 25.000 146.200 ;
        RECT 22.200 142.800 22.600 143.200 ;
        RECT 21.400 138.800 21.800 139.200 ;
        RECT 19.000 135.100 19.400 135.200 ;
        RECT 18.200 134.800 19.400 135.100 ;
        RECT 17.400 106.800 17.800 107.200 ;
        RECT 14.200 73.800 14.600 74.200 ;
        RECT 17.400 73.200 17.700 106.800 ;
        RECT 18.200 81.200 18.500 134.800 ;
        RECT 21.400 103.800 21.800 104.200 ;
        RECT 18.200 80.800 18.600 81.200 ;
        RECT 18.200 73.800 18.600 74.200 ;
        RECT 17.400 72.800 17.800 73.200 ;
        RECT 18.200 67.200 18.500 73.800 ;
        RECT 18.200 66.800 18.600 67.200 ;
        RECT 14.200 66.100 14.600 66.200 ;
        RECT 13.400 65.800 14.600 66.100 ;
        RECT 12.600 50.800 13.000 51.200 ;
        RECT 12.600 46.200 12.900 50.800 ;
        RECT 12.600 45.800 13.000 46.200 ;
        RECT 15.800 36.800 16.200 37.200 ;
        RECT 15.800 36.100 16.100 36.800 ;
        RECT 16.600 36.100 17.000 36.200 ;
        RECT 15.800 35.800 17.000 36.100 ;
        RECT 18.200 35.200 18.500 66.800 ;
        RECT 21.400 37.200 21.700 103.800 ;
        RECT 22.200 96.200 22.500 142.800 ;
        RECT 25.400 108.200 25.700 147.800 ;
        RECT 39.000 134.200 39.300 149.800 ;
        RECT 39.000 133.800 39.400 134.200 ;
        RECT 39.800 131.800 40.200 132.200 ;
        RECT 34.200 125.800 34.600 126.200 ;
        RECT 25.400 107.800 25.800 108.200 ;
        RECT 31.000 107.800 31.400 108.200 ;
        RECT 22.200 95.800 22.600 96.200 ;
        RECT 22.200 48.200 22.500 95.800 ;
        RECT 31.000 92.200 31.300 107.800 ;
        RECT 31.800 105.800 32.200 106.200 ;
        RECT 31.800 105.200 32.100 105.800 ;
        RECT 31.800 104.800 32.200 105.200 ;
        RECT 31.000 91.800 31.400 92.200 ;
        RECT 32.600 88.800 33.000 89.200 ;
        RECT 32.600 72.200 32.900 88.800 ;
        RECT 32.600 71.800 33.000 72.200 ;
        RECT 28.600 70.800 29.000 71.200 ;
        RECT 28.600 66.200 28.900 70.800 ;
        RECT 28.600 65.800 29.000 66.200 ;
        RECT 26.200 58.800 26.600 59.200 ;
        RECT 22.200 47.800 22.600 48.200 ;
        RECT 21.400 36.800 21.800 37.200 ;
        RECT 17.400 34.800 17.800 35.200 ;
        RECT 18.200 34.800 18.600 35.200 ;
        RECT 17.400 26.200 17.700 34.800 ;
        RECT 17.400 25.800 17.800 26.200 ;
        RECT 18.200 15.200 18.500 34.800 ;
        RECT 18.200 14.800 18.600 15.200 ;
        RECT 26.200 12.200 26.500 58.800 ;
        RECT 34.200 57.100 34.500 125.800 ;
        RECT 37.400 123.800 37.800 124.200 ;
        RECT 37.400 91.200 37.700 123.800 ;
        RECT 39.800 108.200 40.100 131.800 ;
        RECT 41.400 130.800 41.800 131.200 ;
        RECT 43.800 130.800 44.200 131.200 ;
        RECT 40.600 127.800 41.000 128.200 ;
        RECT 39.800 107.800 40.200 108.200 ;
        RECT 39.800 96.200 40.100 107.800 ;
        RECT 40.600 99.200 40.900 127.800 ;
        RECT 41.400 109.200 41.700 130.800 ;
        RECT 43.800 129.200 44.100 130.800 ;
        RECT 43.800 128.800 44.200 129.200 ;
        RECT 43.800 123.800 44.200 124.200 ;
        RECT 42.200 114.800 42.600 115.200 ;
        RECT 41.400 108.800 41.800 109.200 ;
        RECT 41.400 107.800 41.800 108.200 ;
        RECT 41.400 106.200 41.700 107.800 ;
        RECT 42.200 106.200 42.500 114.800 ;
        RECT 43.000 106.800 43.400 107.200 ;
        RECT 43.000 106.200 43.300 106.800 ;
        RECT 41.400 105.800 41.800 106.200 ;
        RECT 42.200 105.800 42.600 106.200 ;
        RECT 43.000 105.800 43.400 106.200 ;
        RECT 43.800 104.200 44.100 123.800 ;
        RECT 43.800 103.800 44.200 104.200 ;
        RECT 40.600 98.800 41.000 99.200 ;
        RECT 39.800 95.800 40.200 96.200 ;
        RECT 37.400 90.800 37.800 91.200 ;
        RECT 35.000 57.100 35.400 57.200 ;
        RECT 34.200 56.800 35.400 57.100 ;
        RECT 34.200 55.800 34.600 56.200 ;
        RECT 31.800 47.800 32.200 48.200 ;
        RECT 28.600 36.800 29.000 37.200 ;
        RECT 26.200 11.800 26.600 12.200 ;
        RECT 28.600 9.200 28.900 36.800 ;
        RECT 29.400 34.800 29.800 35.200 ;
        RECT 29.400 34.200 29.700 34.800 ;
        RECT 29.400 33.800 29.800 34.200 ;
        RECT 29.400 31.800 29.800 32.200 ;
        RECT 28.600 8.800 29.000 9.200 ;
        RECT 29.400 8.200 29.700 31.800 ;
        RECT 31.800 18.200 32.100 47.800 ;
        RECT 34.200 29.100 34.500 55.800 ;
        RECT 39.800 37.200 40.100 95.800 ;
        RECT 40.600 92.800 41.000 93.200 ;
        RECT 40.600 56.200 40.900 92.800 ;
        RECT 44.600 87.200 44.900 153.800 ;
        RECT 48.600 129.200 48.900 169.800 ;
        RECT 106.200 167.800 106.600 168.200 ;
        RECT 66.200 164.800 66.600 165.200 ;
        RECT 63.000 157.800 63.400 158.200 ;
        RECT 61.400 150.800 61.800 151.200 ;
        RECT 54.200 145.800 54.600 146.200 ;
        RECT 52.600 133.800 53.000 134.200 ;
        RECT 48.600 128.800 49.000 129.200 ;
        RECT 49.400 129.100 49.800 129.200 ;
        RECT 50.200 129.100 50.600 129.200 ;
        RECT 49.400 128.800 50.600 129.100 ;
        RECT 47.000 126.800 47.400 127.200 ;
        RECT 47.000 126.200 47.300 126.800 ;
        RECT 47.000 125.800 47.400 126.200 ;
        RECT 48.600 110.800 49.000 111.200 ;
        RECT 47.000 95.800 47.400 96.200 ;
        RECT 46.200 93.800 46.600 94.200 ;
        RECT 44.600 86.800 45.000 87.200 ;
        RECT 46.200 68.200 46.500 93.800 ;
        RECT 47.000 81.200 47.300 95.800 ;
        RECT 47.800 94.800 48.200 95.200 ;
        RECT 47.800 94.200 48.100 94.800 ;
        RECT 47.800 93.800 48.200 94.200 ;
        RECT 47.000 80.800 47.400 81.200 ;
        RECT 47.000 76.200 47.300 80.800 ;
        RECT 47.000 75.800 47.400 76.200 ;
        RECT 46.200 67.800 46.600 68.200 ;
        RECT 48.600 67.200 48.900 110.800 ;
        RECT 52.600 77.200 52.900 133.800 ;
        RECT 53.400 122.800 53.800 123.200 ;
        RECT 53.400 97.200 53.700 122.800 ;
        RECT 54.200 114.200 54.500 145.800 ;
        RECT 58.200 127.100 58.600 127.200 ;
        RECT 59.000 127.100 59.400 127.200 ;
        RECT 58.200 126.800 59.400 127.100 ;
        RECT 58.200 116.800 58.600 117.200 ;
        RECT 54.200 113.800 54.600 114.200 ;
        RECT 54.200 106.800 54.600 107.200 ;
        RECT 57.400 106.800 57.800 107.200 ;
        RECT 53.400 96.800 53.800 97.200 ;
        RECT 52.600 76.800 53.000 77.200 ;
        RECT 49.400 76.100 49.800 76.200 ;
        RECT 50.200 76.100 50.600 76.200 ;
        RECT 49.400 75.800 50.600 76.100 ;
        RECT 48.600 66.800 49.000 67.200 ;
        RECT 51.800 66.800 52.200 67.200 ;
        RECT 40.600 55.800 41.000 56.200 ;
        RECT 49.400 46.800 49.800 47.200 ;
        RECT 49.400 45.200 49.700 46.800 ;
        RECT 49.400 44.800 49.800 45.200 ;
        RECT 51.800 44.200 52.100 66.800 ;
        RECT 51.800 43.800 52.200 44.200 ;
        RECT 43.800 41.800 44.200 42.200 ;
        RECT 39.800 36.800 40.200 37.200 ;
        RECT 37.400 36.100 37.800 36.200 ;
        RECT 38.200 36.100 38.600 36.200 ;
        RECT 37.400 35.800 38.600 36.100 ;
        RECT 39.800 35.100 40.200 35.200 ;
        RECT 40.600 35.100 41.000 35.200 ;
        RECT 39.800 34.800 41.000 35.100 ;
        RECT 43.800 33.200 44.100 41.800 ;
        RECT 48.600 34.100 49.000 34.200 ;
        RECT 49.400 34.100 49.800 34.200 ;
        RECT 48.600 33.800 49.800 34.100 ;
        RECT 43.800 32.800 44.200 33.200 ;
        RECT 50.200 29.800 50.600 30.200 ;
        RECT 35.000 29.100 35.400 29.200 ;
        RECT 34.200 28.800 35.400 29.100 ;
        RECT 50.200 25.200 50.500 29.800 ;
        RECT 54.200 26.200 54.500 106.800 ;
        RECT 55.000 74.800 55.400 75.200 ;
        RECT 55.000 65.200 55.300 74.800 ;
        RECT 56.600 72.800 57.000 73.200 ;
        RECT 56.600 70.200 56.900 72.800 ;
        RECT 56.600 69.800 57.000 70.200 ;
        RECT 57.400 69.200 57.700 106.800 ;
        RECT 58.200 83.200 58.500 116.800 ;
        RECT 59.000 94.100 59.400 94.200 ;
        RECT 59.800 94.100 60.200 94.200 ;
        RECT 59.000 93.800 60.200 94.100 ;
        RECT 60.600 88.800 61.000 89.200 ;
        RECT 60.600 84.200 60.900 88.800 ;
        RECT 60.600 83.800 61.000 84.200 ;
        RECT 58.200 82.800 58.600 83.200 ;
        RECT 57.400 68.800 57.800 69.200 ;
        RECT 56.600 65.800 57.000 66.200 ;
        RECT 55.000 64.800 55.400 65.200 ;
        RECT 56.600 44.200 56.900 65.800 ;
        RECT 58.200 56.200 58.500 82.800 ;
        RECT 61.400 82.200 61.700 150.800 ;
        RECT 62.200 148.800 62.600 149.200 ;
        RECT 62.200 99.200 62.500 148.800 ;
        RECT 63.000 148.200 63.300 157.800 ;
        RECT 63.000 147.800 63.400 148.200 ;
        RECT 66.200 135.200 66.500 164.800 ;
        RECT 71.800 163.800 72.200 164.200 ;
        RECT 67.800 141.800 68.200 142.200 ;
        RECT 66.200 134.800 66.600 135.200 ;
        RECT 67.000 131.800 67.400 132.200 ;
        RECT 66.200 128.800 66.600 129.200 ;
        RECT 66.200 127.200 66.500 128.800 ;
        RECT 66.200 126.800 66.600 127.200 ;
        RECT 64.600 117.800 65.000 118.200 ;
        RECT 64.600 108.200 64.900 117.800 ;
        RECT 65.400 115.800 65.800 116.200 ;
        RECT 64.600 107.800 65.000 108.200 ;
        RECT 62.200 98.800 62.600 99.200 ;
        RECT 64.600 94.800 65.000 95.200 ;
        RECT 63.800 93.800 64.200 94.200 ;
        RECT 63.800 93.200 64.100 93.800 ;
        RECT 63.800 92.800 64.200 93.200 ;
        RECT 62.200 82.800 62.600 83.200 ;
        RECT 61.400 81.800 61.800 82.200 ;
        RECT 59.000 74.800 59.400 75.200 ;
        RECT 58.200 55.800 58.600 56.200 ;
        RECT 59.000 55.200 59.300 74.800 ;
        RECT 59.000 54.800 59.400 55.200 ;
        RECT 59.800 53.800 60.200 54.200 ;
        RECT 59.800 51.200 60.100 53.800 ;
        RECT 59.800 50.800 60.200 51.200 ;
        RECT 56.600 43.800 57.000 44.200 ;
        RECT 62.200 40.200 62.500 82.800 ;
        RECT 63.000 67.100 63.400 67.200 ;
        RECT 63.800 67.100 64.200 67.200 ;
        RECT 63.000 66.800 64.200 67.100 ;
        RECT 63.000 54.100 63.400 54.200 ;
        RECT 63.800 54.100 64.200 54.200 ;
        RECT 63.000 53.800 64.200 54.100 ;
        RECT 63.000 41.800 63.400 42.200 ;
        RECT 62.200 39.800 62.600 40.200 ;
        RECT 61.400 35.800 61.800 36.200 ;
        RECT 61.400 34.200 61.700 35.800 ;
        RECT 61.400 33.800 61.800 34.200 ;
        RECT 63.000 27.200 63.300 41.800 ;
        RECT 64.600 41.200 64.900 94.800 ;
        RECT 65.400 89.200 65.700 115.800 ;
        RECT 67.000 107.200 67.300 131.800 ;
        RECT 67.800 113.200 68.100 141.800 ;
        RECT 67.800 112.800 68.200 113.200 ;
        RECT 71.000 110.100 71.400 110.200 ;
        RECT 71.800 110.100 72.100 163.800 ;
        RECT 73.400 162.800 73.800 163.200 ;
        RECT 71.000 109.800 72.100 110.100 ;
        RECT 72.600 109.800 73.000 110.200 ;
        RECT 72.600 108.200 72.900 109.800 ;
        RECT 68.600 108.100 69.000 108.200 ;
        RECT 68.600 107.800 69.700 108.100 ;
        RECT 72.600 107.800 73.000 108.200 ;
        RECT 67.000 106.800 67.400 107.200 ;
        RECT 68.600 105.800 69.000 106.200 ;
        RECT 68.600 101.200 68.900 105.800 ;
        RECT 69.400 105.200 69.700 107.800 ;
        RECT 69.400 104.800 69.800 105.200 ;
        RECT 68.600 100.800 69.000 101.200 ;
        RECT 72.600 96.800 73.000 97.200 ;
        RECT 65.400 88.800 65.800 89.200 ;
        RECT 70.200 88.800 70.600 89.200 ;
        RECT 65.400 87.800 65.800 88.200 ;
        RECT 64.600 40.800 65.000 41.200 ;
        RECT 64.600 35.200 64.900 40.800 ;
        RECT 64.600 34.800 65.000 35.200 ;
        RECT 63.000 26.800 63.400 27.200 ;
        RECT 54.200 25.800 54.600 26.200 ;
        RECT 55.000 26.100 55.400 26.200 ;
        RECT 55.800 26.100 56.200 26.200 ;
        RECT 55.000 25.800 56.200 26.100 ;
        RECT 50.200 24.800 50.600 25.200 ;
        RECT 60.600 25.100 61.000 25.200 ;
        RECT 61.400 25.100 61.800 25.200 ;
        RECT 60.600 24.800 61.800 25.100 ;
        RECT 31.800 17.800 32.200 18.200 ;
        RECT 65.400 17.200 65.700 87.800 ;
        RECT 68.600 84.800 69.000 85.200 ;
        RECT 67.000 74.100 67.400 74.200 ;
        RECT 67.000 73.800 68.100 74.100 ;
        RECT 67.800 53.200 68.100 73.800 ;
        RECT 68.600 59.200 68.900 84.800 ;
        RECT 69.400 77.800 69.800 78.200 ;
        RECT 69.400 72.200 69.700 77.800 ;
        RECT 69.400 71.800 69.800 72.200 ;
        RECT 70.200 66.200 70.500 88.800 ;
        RECT 72.600 77.200 72.900 96.800 ;
        RECT 73.400 95.200 73.700 162.800 ;
        RECT 77.400 159.800 77.800 160.200 ;
        RECT 75.000 149.800 75.400 150.200 ;
        RECT 74.200 96.800 74.600 97.200 ;
        RECT 73.400 94.800 73.800 95.200 ;
        RECT 72.600 76.800 73.000 77.200 ;
        RECT 71.000 76.100 71.400 76.200 ;
        RECT 71.800 76.100 72.200 76.200 ;
        RECT 71.000 75.800 72.200 76.100 ;
        RECT 74.200 75.200 74.500 96.800 ;
        RECT 75.000 86.200 75.300 149.800 ;
        RECT 75.800 131.100 76.200 131.200 ;
        RECT 75.800 130.800 76.900 131.100 ;
        RECT 76.600 122.200 76.900 130.800 ;
        RECT 76.600 121.800 77.000 122.200 ;
        RECT 76.600 99.800 77.000 100.200 ;
        RECT 75.800 97.800 76.200 98.200 ;
        RECT 75.800 95.200 76.100 97.800 ;
        RECT 75.800 94.800 76.200 95.200 ;
        RECT 75.800 90.800 76.200 91.200 ;
        RECT 75.000 85.800 75.400 86.200 ;
        RECT 75.000 75.800 75.400 76.200 ;
        RECT 75.000 75.200 75.300 75.800 ;
        RECT 71.800 74.800 72.200 75.200 ;
        RECT 72.600 74.800 73.000 75.200 ;
        RECT 74.200 74.800 74.600 75.200 ;
        RECT 75.000 74.800 75.400 75.200 ;
        RECT 71.800 73.200 72.100 74.800 ;
        RECT 71.800 72.800 72.200 73.200 ;
        RECT 70.200 65.800 70.600 66.200 ;
        RECT 68.600 58.800 69.000 59.200 ;
        RECT 70.200 53.200 70.500 65.800 ;
        RECT 67.800 52.800 68.200 53.200 ;
        RECT 70.200 52.800 70.600 53.200 ;
        RECT 70.200 35.200 70.500 52.800 ;
        RECT 72.600 50.200 72.900 74.800 ;
        RECT 73.400 74.100 73.800 74.200 ;
        RECT 74.200 74.100 74.600 74.200 ;
        RECT 73.400 73.800 74.600 74.100 ;
        RECT 75.000 73.800 75.400 74.200 ;
        RECT 72.600 49.800 73.000 50.200 ;
        RECT 75.000 37.200 75.300 73.800 ;
        RECT 75.800 70.200 76.100 90.800 ;
        RECT 76.600 75.200 76.900 99.800 ;
        RECT 77.400 79.200 77.700 159.800 ;
        RECT 84.600 158.800 85.000 159.200 ;
        RECT 84.600 148.200 84.900 158.800 ;
        RECT 106.200 155.200 106.500 167.800 ;
        RECT 111.800 155.200 112.100 171.800 ;
        RECT 190.200 167.200 190.500 171.800 ;
        RECT 155.000 166.800 155.400 167.200 ;
        RECT 190.200 166.800 190.600 167.200 ;
        RECT 112.600 165.800 113.000 166.200 ;
        RECT 106.200 154.800 106.600 155.200 ;
        RECT 111.800 154.800 112.200 155.200 ;
        RECT 84.600 147.800 85.000 148.200 ;
        RECT 105.400 144.800 105.800 145.200 ;
        RECT 100.600 142.800 101.000 143.200 ;
        RECT 92.600 140.800 93.000 141.200 ;
        RECT 91.800 135.800 92.200 136.200 ;
        RECT 80.600 132.800 81.000 133.200 ;
        RECT 80.600 102.200 80.900 132.800 ;
        RECT 81.400 132.100 81.800 132.200 ;
        RECT 82.200 132.100 82.600 132.200 ;
        RECT 81.400 131.800 82.600 132.100 ;
        RECT 89.400 128.800 89.800 129.200 ;
        RECT 89.400 128.200 89.700 128.800 ;
        RECT 83.000 128.100 83.400 128.200 ;
        RECT 83.800 128.100 84.200 128.200 ;
        RECT 83.000 127.800 84.200 128.100 ;
        RECT 84.600 127.800 85.000 128.200 ;
        RECT 86.200 128.100 86.600 128.200 ;
        RECT 87.000 128.100 87.400 128.200 ;
        RECT 86.200 127.800 87.400 128.100 ;
        RECT 89.400 127.800 89.800 128.200 ;
        RECT 81.400 120.800 81.800 121.200 ;
        RECT 80.600 101.800 81.000 102.200 ;
        RECT 79.800 93.800 80.200 94.200 ;
        RECT 78.200 85.800 78.600 86.200 ;
        RECT 78.200 85.200 78.500 85.800 ;
        RECT 78.200 84.800 78.600 85.200 ;
        RECT 79.000 84.800 79.400 85.200 ;
        RECT 77.400 78.800 77.800 79.200 ;
        RECT 76.600 74.800 77.000 75.200 ;
        RECT 77.400 74.100 77.800 74.200 ;
        RECT 78.200 74.100 78.600 74.200 ;
        RECT 77.400 73.800 78.600 74.100 ;
        RECT 77.400 73.100 77.800 73.200 ;
        RECT 78.200 73.100 78.600 73.200 ;
        RECT 77.400 72.800 78.600 73.100 ;
        RECT 77.400 71.800 77.800 72.200 ;
        RECT 75.800 69.800 76.200 70.200 ;
        RECT 75.000 36.800 75.400 37.200 ;
        RECT 70.200 34.800 70.600 35.200 ;
        RECT 71.000 34.800 71.400 35.200 ;
        RECT 70.200 30.200 70.500 34.800 ;
        RECT 71.000 33.200 71.300 34.800 ;
        RECT 71.800 33.800 72.200 34.200 ;
        RECT 71.000 32.800 71.400 33.200 ;
        RECT 70.200 29.800 70.600 30.200 ;
        RECT 65.400 16.800 65.800 17.200 ;
        RECT 71.800 14.200 72.100 33.800 ;
        RECT 77.400 32.200 77.700 71.800 ;
        RECT 79.000 58.200 79.300 84.800 ;
        RECT 79.000 57.800 79.400 58.200 ;
        RECT 77.400 31.800 77.800 32.200 ;
        RECT 72.600 26.800 73.000 27.200 ;
        RECT 72.600 26.200 72.900 26.800 ;
        RECT 72.600 25.800 73.000 26.200 ;
        RECT 76.600 26.100 77.000 26.200 ;
        RECT 77.400 26.100 77.800 26.200 ;
        RECT 76.600 25.800 77.800 26.100 ;
        RECT 79.800 22.200 80.100 93.800 ;
        RECT 80.600 91.800 81.000 92.200 ;
        RECT 80.600 36.200 80.900 91.800 ;
        RECT 81.400 66.200 81.700 120.800 ;
        RECT 83.000 94.800 83.400 95.200 ;
        RECT 82.200 93.800 82.600 94.200 ;
        RECT 82.200 86.200 82.500 93.800 ;
        RECT 82.200 85.800 82.600 86.200 ;
        RECT 83.000 81.200 83.300 94.800 ;
        RECT 84.600 89.200 84.900 127.800 ;
        RECT 86.200 117.800 86.600 118.200 ;
        RECT 85.400 104.800 85.800 105.200 ;
        RECT 85.400 93.200 85.700 104.800 ;
        RECT 86.200 98.200 86.500 117.800 ;
        RECT 89.400 100.800 89.800 101.200 ;
        RECT 87.000 98.800 87.400 99.200 ;
        RECT 86.200 97.800 86.600 98.200 ;
        RECT 85.400 92.800 85.800 93.200 ;
        RECT 83.800 88.800 84.200 89.200 ;
        RECT 84.600 88.800 85.000 89.200 ;
        RECT 83.000 80.800 83.400 81.200 ;
        RECT 82.200 74.100 82.600 74.200 ;
        RECT 83.000 74.100 83.400 74.200 ;
        RECT 82.200 73.800 83.400 74.100 ;
        RECT 81.400 65.800 81.800 66.200 ;
        RECT 83.800 62.200 84.100 88.800 ;
        RECT 87.000 86.200 87.300 98.800 ;
        RECT 87.000 85.800 87.400 86.200 ;
        RECT 84.600 74.800 85.000 75.200 ;
        RECT 84.600 73.200 84.900 74.800 ;
        RECT 84.600 72.800 85.000 73.200 ;
        RECT 84.600 67.100 85.000 67.200 ;
        RECT 85.400 67.100 85.800 67.200 ;
        RECT 84.600 66.800 85.800 67.100 ;
        RECT 83.800 61.800 84.200 62.200 ;
        RECT 87.000 52.200 87.300 85.800 ;
        RECT 87.800 75.100 88.200 75.200 ;
        RECT 88.600 75.100 89.000 75.200 ;
        RECT 87.800 74.800 89.000 75.100 ;
        RECT 88.600 63.800 89.000 64.200 ;
        RECT 87.800 55.800 88.200 56.200 ;
        RECT 87.000 51.800 87.400 52.200 ;
        RECT 87.000 49.200 87.300 51.800 ;
        RECT 87.000 48.800 87.400 49.200 ;
        RECT 86.200 45.800 86.600 46.200 ;
        RECT 84.600 41.800 85.000 42.200 ;
        RECT 81.400 37.100 81.800 37.200 ;
        RECT 82.200 37.100 82.600 37.200 ;
        RECT 81.400 36.800 82.600 37.100 ;
        RECT 80.600 35.800 81.000 36.200 ;
        RECT 81.400 28.100 81.800 28.200 ;
        RECT 82.200 28.100 82.600 28.200 ;
        RECT 81.400 27.800 82.600 28.100 ;
        RECT 79.800 21.800 80.200 22.200 ;
        RECT 71.800 13.800 72.200 14.200 ;
        RECT 84.600 11.200 84.900 41.800 ;
        RECT 84.600 10.800 85.000 11.200 ;
        RECT 86.200 10.200 86.500 45.800 ;
        RECT 87.800 17.200 88.100 55.800 ;
        RECT 88.600 46.200 88.900 63.800 ;
        RECT 88.600 45.800 89.000 46.200 ;
        RECT 89.400 45.200 89.700 100.800 ;
        RECT 91.800 98.100 92.100 135.800 ;
        RECT 92.600 116.200 92.900 140.800 ;
        RECT 95.800 135.800 96.200 136.200 ;
        RECT 92.600 115.800 93.000 116.200 ;
        RECT 92.600 107.100 93.000 107.200 ;
        RECT 93.400 107.100 93.800 107.200 ;
        RECT 92.600 106.800 93.800 107.100 ;
        RECT 95.800 106.200 96.100 135.800 ;
        RECT 99.000 132.100 99.400 132.200 ;
        RECT 99.800 132.100 100.200 132.200 ;
        RECT 99.000 131.800 100.200 132.100 ;
        RECT 99.800 114.800 100.200 115.200 ;
        RECT 95.800 105.800 96.200 106.200 ;
        RECT 92.600 98.100 93.000 98.200 ;
        RECT 91.800 97.800 93.000 98.100 ;
        RECT 99.800 94.200 100.100 114.800 ;
        RECT 93.400 93.800 93.800 94.200 ;
        RECT 99.800 93.800 100.200 94.200 ;
        RECT 90.200 92.800 90.600 93.200 ;
        RECT 90.200 72.200 90.500 92.800 ;
        RECT 91.800 74.100 92.200 74.200 ;
        RECT 91.000 73.800 92.200 74.100 ;
        RECT 91.000 73.200 91.300 73.800 ;
        RECT 91.000 72.800 91.400 73.200 ;
        RECT 90.200 71.800 90.600 72.200 ;
        RECT 92.600 66.800 93.000 67.200 ;
        RECT 92.600 66.200 92.900 66.800 ;
        RECT 92.600 65.800 93.000 66.200 ;
        RECT 93.400 64.200 93.700 93.800 ;
        RECT 99.000 87.100 99.400 87.200 ;
        RECT 99.800 87.100 100.200 87.200 ;
        RECT 99.000 86.800 100.200 87.100 ;
        RECT 100.600 85.200 100.900 142.800 ;
        RECT 103.800 126.800 104.200 127.200 ;
        RECT 100.600 84.800 101.000 85.200 ;
        RECT 95.000 81.800 95.400 82.200 ;
        RECT 93.400 63.800 93.800 64.200 ;
        RECT 90.200 61.800 90.600 62.200 ;
        RECT 90.200 50.200 90.500 61.800 ;
        RECT 90.200 49.800 90.600 50.200 ;
        RECT 91.000 49.100 91.400 49.200 ;
        RECT 91.800 49.100 92.200 49.200 ;
        RECT 91.000 48.800 92.200 49.100 ;
        RECT 89.400 44.800 89.800 45.200 ;
        RECT 90.200 42.800 90.600 43.200 ;
        RECT 90.200 27.200 90.500 42.800 ;
        RECT 95.000 35.200 95.300 81.800 ;
        RECT 95.800 79.800 96.200 80.200 ;
        RECT 95.800 65.200 96.100 79.800 ;
        RECT 100.600 77.800 101.000 78.200 ;
        RECT 99.000 76.800 99.400 77.200 ;
        RECT 98.200 69.100 98.600 69.200 ;
        RECT 99.000 69.100 99.300 76.800 ;
        RECT 98.200 68.800 99.300 69.100 ;
        RECT 99.800 68.800 100.200 69.200 ;
        RECT 99.800 67.200 100.100 68.800 ;
        RECT 99.800 66.800 100.200 67.200 ;
        RECT 95.800 64.800 96.200 65.200 ;
        RECT 95.000 34.800 95.400 35.200 ;
        RECT 91.800 27.800 92.200 28.200 ;
        RECT 93.400 28.100 93.800 28.200 ;
        RECT 94.200 28.100 94.600 28.200 ;
        RECT 93.400 27.800 94.600 28.100 ;
        RECT 91.800 27.200 92.100 27.800 ;
        RECT 95.000 27.200 95.300 34.800 ;
        RECT 95.800 34.200 96.100 64.800 ;
        RECT 99.800 52.800 100.200 53.200 ;
        RECT 97.400 46.800 97.800 47.200 ;
        RECT 96.600 45.800 97.000 46.200 ;
        RECT 97.400 46.100 97.700 46.800 ;
        RECT 98.200 46.100 98.600 46.200 ;
        RECT 97.400 45.800 98.600 46.100 ;
        RECT 95.800 33.800 96.200 34.200 ;
        RECT 95.800 27.200 96.100 33.800 ;
        RECT 96.600 31.200 96.900 45.800 ;
        RECT 99.800 45.200 100.100 52.800 ;
        RECT 100.600 46.200 100.900 77.800 ;
        RECT 103.800 59.200 104.100 126.800 ;
        RECT 105.400 115.200 105.700 144.800 ;
        RECT 107.800 138.800 108.200 139.200 ;
        RECT 106.200 126.800 106.600 127.200 ;
        RECT 106.200 126.200 106.500 126.800 ;
        RECT 106.200 125.800 106.600 126.200 ;
        RECT 105.400 114.800 105.800 115.200 ;
        RECT 104.600 100.800 105.000 101.200 ;
        RECT 104.600 91.200 104.900 100.800 ;
        RECT 104.600 90.800 105.000 91.200 ;
        RECT 104.600 88.800 105.000 89.200 ;
        RECT 103.800 58.800 104.200 59.200 ;
        RECT 104.600 52.200 104.900 88.800 ;
        RECT 105.400 87.100 105.800 87.200 ;
        RECT 106.200 87.100 106.600 87.200 ;
        RECT 105.400 86.800 106.600 87.100 ;
        RECT 107.000 75.800 107.400 76.200 ;
        RECT 105.400 74.800 105.800 75.200 ;
        RECT 106.200 74.800 106.600 75.200 ;
        RECT 104.600 51.800 105.000 52.200 ;
        RECT 104.600 49.800 105.000 50.200 ;
        RECT 104.600 47.200 104.900 49.800 ;
        RECT 105.400 47.200 105.700 74.800 ;
        RECT 106.200 74.200 106.500 74.800 ;
        RECT 106.200 73.800 106.600 74.200 ;
        RECT 103.800 46.800 104.200 47.200 ;
        RECT 104.600 46.800 105.000 47.200 ;
        RECT 105.400 46.800 105.800 47.200 ;
        RECT 106.200 46.800 106.600 47.200 ;
        RECT 100.600 45.800 101.000 46.200 ;
        RECT 99.800 44.800 100.200 45.200 ;
        RECT 98.200 36.800 98.600 37.200 ;
        RECT 98.200 35.200 98.500 36.800 ;
        RECT 98.200 34.800 98.600 35.200 ;
        RECT 96.600 30.800 97.000 31.200 ;
        RECT 90.200 26.800 90.600 27.200 ;
        RECT 91.800 26.800 92.200 27.200 ;
        RECT 92.600 26.800 93.000 27.200 ;
        RECT 95.000 26.800 95.400 27.200 ;
        RECT 95.800 26.800 96.200 27.200 ;
        RECT 92.600 26.200 92.900 26.800 ;
        RECT 98.200 26.200 98.500 34.800 ;
        RECT 100.600 29.800 101.000 30.200 ;
        RECT 92.600 25.800 93.000 26.200 ;
        RECT 98.200 25.800 98.600 26.200 ;
        RECT 99.800 26.100 100.200 26.200 ;
        RECT 100.600 26.100 100.900 29.800 ;
        RECT 99.800 25.800 100.900 26.100 ;
        RECT 103.800 26.200 104.100 46.800 ;
        RECT 104.600 45.800 105.000 46.200 ;
        RECT 104.600 32.200 104.900 45.800 ;
        RECT 106.200 40.200 106.500 46.800 ;
        RECT 106.200 39.800 106.600 40.200 ;
        RECT 105.400 34.100 105.800 34.200 ;
        RECT 106.200 34.100 106.600 34.200 ;
        RECT 105.400 33.800 106.600 34.100 ;
        RECT 104.600 31.800 105.000 32.200 ;
        RECT 104.600 28.800 105.000 29.200 ;
        RECT 104.600 28.200 104.900 28.800 ;
        RECT 104.600 27.800 105.000 28.200 ;
        RECT 103.800 25.800 104.200 26.200 ;
        RECT 103.800 24.200 104.100 25.800 ;
        RECT 103.800 23.800 104.200 24.200 ;
        RECT 88.600 18.800 89.000 19.200 ;
        RECT 88.600 17.200 88.900 18.800 ;
        RECT 87.800 16.800 88.200 17.200 ;
        RECT 88.600 16.800 89.000 17.200 ;
        RECT 107.000 16.200 107.300 75.800 ;
        RECT 107.800 50.200 108.100 138.800 ;
        RECT 109.400 128.800 109.800 129.200 ;
        RECT 109.400 128.200 109.700 128.800 ;
        RECT 109.400 127.800 109.800 128.200 ;
        RECT 112.600 104.200 112.900 165.800 ;
        RECT 123.000 161.800 123.400 162.200 ;
        RECT 120.600 144.800 121.000 145.200 ;
        RECT 115.800 141.800 116.200 142.200 ;
        RECT 115.000 130.800 115.400 131.200 ;
        RECT 113.400 123.800 113.800 124.200 ;
        RECT 112.600 103.800 113.000 104.200 ;
        RECT 113.400 103.200 113.700 123.800 ;
        RECT 113.400 102.800 113.800 103.200 ;
        RECT 115.000 89.200 115.300 130.800 ;
        RECT 115.800 128.200 116.100 141.800 ;
        RECT 120.600 136.200 120.900 144.800 ;
        RECT 123.000 143.200 123.300 161.800 ;
        RECT 151.800 153.800 152.200 154.200 ;
        RECT 138.200 152.800 138.600 153.200 ;
        RECT 125.400 149.800 125.800 150.200 ;
        RECT 123.800 146.800 124.200 147.200 ;
        RECT 123.000 142.800 123.400 143.200 ;
        RECT 120.600 135.800 121.000 136.200 ;
        RECT 122.200 135.100 122.600 135.200 ;
        RECT 123.000 135.100 123.400 135.200 ;
        RECT 122.200 134.800 123.400 135.100 ;
        RECT 115.800 127.800 116.200 128.200 ;
        RECT 115.800 113.200 116.100 127.800 ;
        RECT 119.000 115.800 119.400 116.200 ;
        RECT 117.400 114.100 117.800 114.200 ;
        RECT 118.200 114.100 118.600 114.200 ;
        RECT 117.400 113.800 118.600 114.100 ;
        RECT 115.800 112.800 116.200 113.200 ;
        RECT 115.800 92.200 116.100 112.800 ;
        RECT 116.600 102.800 117.000 103.200 ;
        RECT 115.800 91.800 116.200 92.200 ;
        RECT 115.000 88.800 115.400 89.200 ;
        RECT 115.000 76.200 115.300 88.800 ;
        RECT 115.800 78.800 116.200 79.200 ;
        RECT 115.000 75.800 115.400 76.200 ;
        RECT 111.000 72.800 111.400 73.200 ;
        RECT 110.200 56.800 110.600 57.200 ;
        RECT 108.600 50.800 109.000 51.200 ;
        RECT 107.800 49.800 108.200 50.200 ;
        RECT 108.600 48.200 108.900 50.800 ;
        RECT 109.400 49.800 109.800 50.200 ;
        RECT 108.600 47.800 109.000 48.200 ;
        RECT 108.600 46.800 109.000 47.200 ;
        RECT 108.600 44.200 108.900 46.800 ;
        RECT 108.600 43.800 109.000 44.200 ;
        RECT 109.400 40.200 109.700 49.800 ;
        RECT 109.400 39.800 109.800 40.200 ;
        RECT 108.600 37.100 109.000 37.200 ;
        RECT 109.400 37.100 109.800 37.200 ;
        RECT 108.600 36.800 109.800 37.100 ;
        RECT 107.000 15.800 107.400 16.200 ;
        RECT 110.200 13.200 110.500 56.800 ;
        RECT 111.000 17.200 111.300 72.800 ;
        RECT 111.800 53.800 112.200 54.200 ;
        RECT 111.800 27.200 112.100 53.800 ;
        RECT 115.000 51.800 115.400 52.200 ;
        RECT 114.200 51.100 114.600 51.200 ;
        RECT 115.000 51.100 115.300 51.800 ;
        RECT 114.200 50.800 115.300 51.100 ;
        RECT 113.400 48.800 113.800 49.200 ;
        RECT 113.400 47.200 113.700 48.800 ;
        RECT 113.400 46.800 113.800 47.200 ;
        RECT 112.600 37.100 113.000 37.200 ;
        RECT 113.400 37.100 113.800 37.200 ;
        RECT 112.600 36.800 113.800 37.100 ;
        RECT 115.000 30.200 115.300 50.800 ;
        RECT 115.800 45.200 116.100 78.800 ;
        RECT 116.600 72.200 116.900 102.800 ;
        RECT 119.000 79.200 119.300 115.800 ;
        RECT 123.800 106.200 124.100 146.800 ;
        RECT 125.400 136.200 125.700 149.800 ;
        RECT 127.800 142.800 128.200 143.200 ;
        RECT 127.800 139.200 128.100 142.800 ;
        RECT 128.600 140.800 129.000 141.200 ;
        RECT 127.800 138.800 128.200 139.200 ;
        RECT 127.000 136.800 127.400 137.200 ;
        RECT 125.400 135.800 125.800 136.200 ;
        RECT 123.800 105.800 124.200 106.200 ;
        RECT 121.400 103.800 121.800 104.200 ;
        RECT 119.000 78.800 119.400 79.200 ;
        RECT 119.000 77.800 119.400 78.200 ;
        RECT 116.600 71.800 117.000 72.200 ;
        RECT 119.000 68.200 119.300 77.800 ;
        RECT 119.000 67.800 119.400 68.200 ;
        RECT 118.200 58.800 118.600 59.200 ;
        RECT 116.600 56.800 117.000 57.200 ;
        RECT 116.600 46.200 116.900 56.800 ;
        RECT 117.400 53.800 117.800 54.200 ;
        RECT 117.400 52.200 117.700 53.800 ;
        RECT 117.400 51.800 117.800 52.200 ;
        RECT 116.600 45.800 117.000 46.200 ;
        RECT 115.800 44.800 116.200 45.200 ;
        RECT 116.600 33.800 117.000 34.200 ;
        RECT 116.600 33.200 116.900 33.800 ;
        RECT 116.600 32.800 117.000 33.200 ;
        RECT 115.000 29.800 115.400 30.200 ;
        RECT 117.400 27.800 117.800 28.200 ;
        RECT 117.400 27.200 117.700 27.800 ;
        RECT 111.800 26.800 112.200 27.200 ;
        RECT 117.400 26.800 117.800 27.200 ;
        RECT 114.200 25.800 114.600 26.200 ;
        RECT 114.200 20.200 114.500 25.800 ;
        RECT 118.200 25.200 118.500 58.800 ;
        RECT 119.000 54.800 119.400 55.200 ;
        RECT 119.000 41.200 119.300 54.800 ;
        RECT 120.600 53.800 121.000 54.200 ;
        RECT 119.000 40.800 119.400 41.200 ;
        RECT 118.200 24.800 118.600 25.200 ;
        RECT 114.200 19.800 114.600 20.200 ;
        RECT 111.000 16.800 111.400 17.200 ;
        RECT 115.800 17.100 116.200 17.200 ;
        RECT 115.000 16.800 116.200 17.100 ;
        RECT 110.200 12.800 110.600 13.200 ;
        RECT 86.200 9.800 86.600 10.200 ;
        RECT 115.000 9.200 115.300 16.800 ;
        RECT 119.000 14.200 119.300 40.800 ;
        RECT 120.600 34.200 120.900 53.800 ;
        RECT 120.600 33.800 121.000 34.200 ;
        RECT 119.000 13.800 119.400 14.200 ;
        RECT 115.000 8.800 115.400 9.200 ;
        RECT 29.400 7.800 29.800 8.200 ;
        RECT 29.400 6.200 29.700 7.800 ;
        RECT 121.400 7.200 121.700 103.800 ;
        RECT 126.200 96.800 126.600 97.200 ;
        RECT 123.800 73.800 124.200 74.200 ;
        RECT 122.200 71.800 122.600 72.200 ;
        RECT 122.200 25.200 122.500 71.800 ;
        RECT 123.800 63.200 124.100 73.800 ;
        RECT 123.800 62.800 124.200 63.200 ;
        RECT 126.200 62.200 126.500 96.800 ;
        RECT 127.000 65.200 127.300 136.800 ;
        RECT 128.600 134.200 128.900 140.800 ;
        RECT 136.600 135.100 137.000 135.200 ;
        RECT 137.400 135.100 137.800 135.200 ;
        RECT 136.600 134.800 137.800 135.100 ;
        RECT 128.600 133.800 129.000 134.200 ;
        RECT 128.600 111.200 128.900 133.800 ;
        RECT 135.800 131.800 136.200 132.200 ;
        RECT 135.800 130.200 136.100 131.800 ;
        RECT 135.800 129.800 136.200 130.200 ;
        RECT 138.200 115.200 138.500 152.800 ;
        RECT 147.000 140.800 147.400 141.200 ;
        RECT 139.000 126.800 139.400 127.200 ;
        RECT 129.400 114.800 129.800 115.200 ;
        RECT 138.200 114.800 138.600 115.200 ;
        RECT 128.600 110.800 129.000 111.200 ;
        RECT 129.400 108.200 129.700 114.800 ;
        RECT 130.200 114.100 130.600 114.200 ;
        RECT 131.000 114.100 131.400 114.200 ;
        RECT 130.200 113.800 131.400 114.100 ;
        RECT 129.400 107.800 129.800 108.200 ;
        RECT 139.000 95.200 139.300 126.800 ;
        RECT 139.800 125.800 140.200 126.200 ;
        RECT 139.000 94.800 139.400 95.200 ;
        RECT 139.000 87.200 139.300 94.800 ;
        RECT 139.000 86.800 139.400 87.200 ;
        RECT 129.400 74.800 129.800 75.200 ;
        RECT 129.400 73.200 129.700 74.800 ;
        RECT 129.400 72.800 129.800 73.200 ;
        RECT 128.600 67.800 129.000 68.200 ;
        RECT 134.200 68.100 134.600 68.200 ;
        RECT 135.000 68.100 135.400 68.200 ;
        RECT 134.200 67.800 135.400 68.100 ;
        RECT 128.600 67.200 128.900 67.800 ;
        RECT 128.600 66.800 129.000 67.200 ;
        RECT 135.800 65.800 136.200 66.200 ;
        RECT 127.000 64.800 127.400 65.200 ;
        RECT 135.800 62.200 136.100 65.800 ;
        RECT 126.200 61.800 126.600 62.200 ;
        RECT 135.800 61.800 136.200 62.200 ;
        RECT 139.000 61.200 139.300 86.800 ;
        RECT 139.800 77.100 140.100 125.800 ;
        RECT 145.400 115.800 145.800 116.200 ;
        RECT 145.400 95.200 145.700 115.800 ;
        RECT 146.200 112.800 146.600 113.200 ;
        RECT 146.200 95.200 146.500 112.800 ;
        RECT 147.000 107.200 147.300 140.800 ;
        RECT 151.800 134.200 152.100 153.800 ;
        RECT 155.000 146.200 155.300 166.800 ;
        RECT 169.400 159.800 169.800 160.200 ;
        RECT 169.400 149.200 169.700 159.800 ;
        RECT 190.200 153.800 190.600 154.200 ;
        RECT 175.000 152.800 175.400 153.200 ;
        RECT 169.400 148.800 169.800 149.200 ;
        RECT 174.200 146.800 174.600 147.200 ;
        RECT 155.000 145.800 155.400 146.200 ;
        RECT 171.000 144.800 171.400 145.200 ;
        RECT 161.400 141.800 161.800 142.200 ;
        RECT 151.800 133.800 152.200 134.200 ;
        RECT 151.800 129.800 152.200 130.200 ;
        RECT 151.000 114.800 151.400 115.200 ;
        RECT 151.000 110.200 151.300 114.800 ;
        RECT 151.000 109.800 151.400 110.200 ;
        RECT 147.000 106.800 147.400 107.200 ;
        RECT 148.600 101.800 149.000 102.200 ;
        RECT 145.400 94.800 145.800 95.200 ;
        RECT 146.200 94.800 146.600 95.200 ;
        RECT 147.800 88.800 148.200 89.200 ;
        RECT 143.800 86.100 144.200 86.200 ;
        RECT 144.600 86.100 145.000 86.200 ;
        RECT 143.800 85.800 145.000 86.100 ;
        RECT 140.600 77.100 141.000 77.200 ;
        RECT 139.800 76.800 141.000 77.100 ;
        RECT 142.200 73.800 142.600 74.200 ;
        RECT 143.800 74.100 144.200 74.200 ;
        RECT 144.600 74.100 145.000 74.200 ;
        RECT 143.800 73.800 145.000 74.100 ;
        RECT 142.200 73.200 142.500 73.800 ;
        RECT 142.200 72.800 142.600 73.200 ;
        RECT 143.800 73.100 144.200 73.200 ;
        RECT 144.600 73.100 145.000 73.200 ;
        RECT 143.800 72.800 145.000 73.100 ;
        RECT 146.200 68.100 146.600 68.200 ;
        RECT 147.000 68.100 147.400 68.200 ;
        RECT 146.200 67.800 147.400 68.100 ;
        RECT 139.000 60.800 139.400 61.200 ;
        RECT 147.800 47.200 148.100 88.800 ;
        RECT 148.600 59.200 148.900 101.800 ;
        RECT 150.200 94.100 150.600 94.200 ;
        RECT 150.200 93.800 151.300 94.100 ;
        RECT 151.000 70.200 151.300 93.800 ;
        RECT 151.000 69.800 151.400 70.200 ;
        RECT 149.400 66.800 149.800 67.200 ;
        RECT 151.800 67.100 152.100 129.800 ;
        RECT 155.000 129.100 155.400 129.200 ;
        RECT 155.800 129.100 156.200 129.200 ;
        RECT 155.000 128.800 156.200 129.100 ;
        RECT 158.200 127.100 158.600 127.200 ;
        RECT 159.000 127.100 159.400 127.200 ;
        RECT 158.200 126.800 159.400 127.100 ;
        RECT 161.400 126.200 161.700 141.800 ;
        RECT 164.600 136.800 165.000 137.200 ;
        RECT 161.400 125.800 161.800 126.200 ;
        RECT 163.000 121.800 163.400 122.200 ;
        RECT 159.800 119.800 160.200 120.200 ;
        RECT 157.400 115.800 157.800 116.200 ;
        RECT 153.400 93.100 153.800 93.200 ;
        RECT 154.200 93.100 154.600 93.200 ;
        RECT 153.400 92.800 154.600 93.100 ;
        RECT 154.200 74.100 154.600 74.200 ;
        RECT 155.000 74.100 155.400 74.200 ;
        RECT 154.200 73.800 155.400 74.100 ;
        RECT 152.600 67.100 153.000 67.200 ;
        RECT 151.800 66.800 153.000 67.100 ;
        RECT 148.600 58.800 149.000 59.200 ;
        RECT 148.600 48.800 149.000 49.200 ;
        RECT 148.600 48.200 148.900 48.800 ;
        RECT 148.600 47.800 149.000 48.200 ;
        RECT 147.800 46.800 148.200 47.200 ;
        RECT 149.400 46.200 149.700 66.800 ;
        RECT 155.000 46.800 155.400 47.200 ;
        RECT 149.400 45.800 149.800 46.200 ;
        RECT 149.400 45.200 149.700 45.800 ;
        RECT 127.000 45.100 127.400 45.200 ;
        RECT 126.200 44.800 127.400 45.100 ;
        RECT 127.800 44.800 128.200 45.200 ;
        RECT 149.400 44.800 149.800 45.200 ;
        RECT 123.800 26.100 124.200 26.200 ;
        RECT 124.600 26.100 125.000 26.200 ;
        RECT 123.800 25.800 125.000 26.100 ;
        RECT 122.200 24.800 122.600 25.200 ;
        RECT 126.200 24.200 126.500 44.800 ;
        RECT 126.200 23.800 126.600 24.200 ;
        RECT 127.800 21.200 128.100 44.800 ;
        RECT 155.000 41.200 155.300 46.800 ;
        RECT 156.600 43.800 157.000 44.200 ;
        RECT 155.000 40.800 155.400 41.200 ;
        RECT 156.600 36.200 156.900 43.800 ;
        RECT 156.600 35.800 157.000 36.200 ;
        RECT 127.800 20.800 128.200 21.200 ;
        RECT 157.400 10.200 157.700 115.800 ;
        RECT 159.000 92.800 159.400 93.200 ;
        RECT 159.000 84.200 159.300 92.800 ;
        RECT 159.800 91.200 160.100 119.800 ;
        RECT 160.600 114.800 161.000 115.200 ;
        RECT 159.800 90.800 160.200 91.200 ;
        RECT 159.800 88.800 160.200 89.200 ;
        RECT 159.800 86.200 160.100 88.800 ;
        RECT 159.800 85.800 160.200 86.200 ;
        RECT 159.000 83.800 159.400 84.200 ;
        RECT 160.600 77.200 160.900 114.800 ;
        RECT 162.200 96.800 162.600 97.200 ;
        RECT 162.200 94.200 162.500 96.800 ;
        RECT 162.200 93.800 162.600 94.200 ;
        RECT 162.200 84.800 162.600 85.200 ;
        RECT 160.600 76.800 161.000 77.200 ;
        RECT 158.200 75.800 158.600 76.200 ;
        RECT 161.400 75.800 161.800 76.200 ;
        RECT 158.200 74.200 158.500 75.800 ;
        RECT 159.800 74.800 160.200 75.200 ;
        RECT 158.200 73.800 158.600 74.200 ;
        RECT 159.800 18.100 160.100 74.800 ;
        RECT 161.400 66.200 161.700 75.800 ;
        RECT 161.400 65.800 161.800 66.200 ;
        RECT 162.200 44.200 162.500 84.800 ;
        RECT 163.000 82.200 163.300 121.800 ;
        RECT 164.600 114.200 164.900 136.800 ;
        RECT 165.400 132.800 165.800 133.200 ;
        RECT 164.600 113.800 165.000 114.200 ;
        RECT 163.800 112.800 164.200 113.200 ;
        RECT 163.000 81.800 163.400 82.200 ;
        RECT 163.800 81.100 164.100 112.800 ;
        RECT 165.400 107.200 165.700 132.800 ;
        RECT 168.600 127.100 169.000 127.200 ;
        RECT 169.400 127.100 169.800 127.200 ;
        RECT 168.600 126.800 169.800 127.100 ;
        RECT 171.000 124.200 171.300 144.800 ;
        RECT 173.400 141.100 173.800 141.200 ;
        RECT 172.600 140.800 173.800 141.100 ;
        RECT 172.600 124.200 172.900 140.800 ;
        RECT 173.400 139.800 173.800 140.200 ;
        RECT 171.000 123.800 171.400 124.200 ;
        RECT 171.800 123.800 172.200 124.200 ;
        RECT 172.600 123.800 173.000 124.200 ;
        RECT 166.200 107.800 166.600 108.200 ;
        RECT 169.400 108.100 169.800 108.200 ;
        RECT 170.200 108.100 170.600 108.200 ;
        RECT 169.400 107.800 170.600 108.100 ;
        RECT 166.200 107.200 166.500 107.800 ;
        RECT 165.400 107.100 165.800 107.200 ;
        RECT 163.000 80.800 164.100 81.100 ;
        RECT 164.600 106.800 165.800 107.100 ;
        RECT 166.200 106.800 166.600 107.200 ;
        RECT 162.200 43.800 162.600 44.200 ;
        RECT 160.600 18.100 161.000 18.200 ;
        RECT 159.800 17.800 161.000 18.100 ;
        RECT 163.000 14.200 163.300 80.800 ;
        RECT 163.800 72.800 164.200 73.200 ;
        RECT 163.800 53.200 164.100 72.800 ;
        RECT 164.600 66.200 164.900 106.800 ;
        RECT 171.800 106.200 172.100 123.800 ;
        RECT 173.400 121.200 173.700 139.800 ;
        RECT 174.200 126.200 174.500 146.800 ;
        RECT 174.200 125.800 174.600 126.200 ;
        RECT 173.400 120.800 173.800 121.200 ;
        RECT 175.000 113.200 175.300 152.800 ;
        RECT 182.200 150.100 182.600 150.200 ;
        RECT 182.200 149.800 183.300 150.100 ;
        RECT 183.000 145.200 183.300 149.800 ;
        RECT 183.800 149.800 184.200 150.200 ;
        RECT 183.000 144.800 183.400 145.200 ;
        RECT 179.000 134.100 179.400 134.200 ;
        RECT 179.800 134.100 180.200 134.200 ;
        RECT 179.000 133.800 180.200 134.100 ;
        RECT 176.600 129.800 177.000 130.200 ;
        RECT 175.800 129.100 176.200 129.200 ;
        RECT 176.600 129.100 176.900 129.800 ;
        RECT 175.800 128.800 176.900 129.100 ;
        RECT 183.800 125.200 184.100 149.800 ;
        RECT 185.400 145.800 185.800 146.200 ;
        RECT 185.400 144.200 185.700 145.800 ;
        RECT 190.200 145.200 190.500 153.800 ;
        RECT 196.600 151.200 196.900 172.800 ;
        RECT 201.400 165.800 201.800 166.200 ;
        RECT 197.400 163.800 197.800 164.200 ;
        RECT 196.600 150.800 197.000 151.200 ;
        RECT 190.200 144.800 190.600 145.200 ;
        RECT 185.400 143.800 185.800 144.200 ;
        RECT 183.800 124.800 184.200 125.200 ;
        RECT 188.600 121.800 189.000 122.200 ;
        RECT 175.000 112.800 175.400 113.200 ;
        RECT 172.600 108.800 173.000 109.200 ;
        RECT 172.600 108.200 172.900 108.800 ;
        RECT 172.600 107.800 173.000 108.200 ;
        RECT 171.800 105.800 172.200 106.200 ;
        RECT 179.800 105.100 180.200 105.200 ;
        RECT 179.800 104.800 180.900 105.100 ;
        RECT 169.400 98.800 169.800 99.200 ;
        RECT 165.400 93.800 165.800 94.200 ;
        RECT 164.600 65.800 165.000 66.200 ;
        RECT 164.600 56.200 164.900 65.800 ;
        RECT 164.600 55.800 165.000 56.200 ;
        RECT 163.800 52.800 164.200 53.200 ;
        RECT 164.600 45.200 164.900 55.800 ;
        RECT 164.600 44.800 165.000 45.200 ;
        RECT 164.600 37.200 164.900 44.800 ;
        RECT 165.400 42.200 165.700 93.800 ;
        RECT 166.200 85.800 166.600 86.200 ;
        RECT 166.200 85.200 166.500 85.800 ;
        RECT 166.200 84.800 166.600 85.200 ;
        RECT 168.600 82.800 169.000 83.200 ;
        RECT 166.200 67.800 166.600 68.200 ;
        RECT 167.800 67.800 168.200 68.200 ;
        RECT 166.200 67.200 166.500 67.800 ;
        RECT 167.800 67.200 168.100 67.800 ;
        RECT 166.200 66.800 166.600 67.200 ;
        RECT 167.800 66.800 168.200 67.200 ;
        RECT 168.600 66.200 168.900 82.800 ;
        RECT 169.400 73.200 169.700 98.800 ;
        RECT 170.200 86.800 170.600 87.200 ;
        RECT 175.800 87.100 176.200 87.200 ;
        RECT 176.600 87.100 177.000 87.200 ;
        RECT 175.800 86.800 177.000 87.100 ;
        RECT 170.200 74.200 170.500 86.800 ;
        RECT 170.200 73.800 170.600 74.200 ;
        RECT 169.400 72.800 169.800 73.200 ;
        RECT 180.600 72.200 180.900 104.800 ;
        RECT 180.600 71.800 181.000 72.200 ;
        RECT 168.600 65.800 169.000 66.200 ;
        RECT 188.600 55.200 188.900 121.800 ;
        RECT 188.600 54.800 189.000 55.200 ;
        RECT 190.200 42.200 190.500 144.800 ;
        RECT 195.800 141.800 196.200 142.200 ;
        RECT 195.800 134.200 196.100 141.800 ;
        RECT 197.400 134.200 197.700 163.800 ;
        RECT 201.400 145.200 201.700 165.800 ;
        RECT 201.400 144.800 201.800 145.200 ;
        RECT 199.800 142.800 200.200 143.200 ;
        RECT 199.800 141.200 200.100 142.800 ;
        RECT 199.800 140.800 200.200 141.200 ;
        RECT 199.000 135.800 199.400 136.200 ;
        RECT 195.800 133.800 196.200 134.200 ;
        RECT 197.400 133.800 197.800 134.200 ;
        RECT 191.000 121.800 191.400 122.200 ;
        RECT 191.000 101.200 191.300 121.800 ;
        RECT 194.200 111.800 194.600 112.200 ;
        RECT 193.400 109.800 193.800 110.200 ;
        RECT 192.600 105.800 193.000 106.200 ;
        RECT 191.000 100.800 191.400 101.200 ;
        RECT 191.000 86.100 191.400 86.200 ;
        RECT 191.800 86.100 192.200 86.200 ;
        RECT 191.000 85.800 192.200 86.100 ;
        RECT 192.600 50.200 192.900 105.800 ;
        RECT 193.400 73.200 193.700 109.800 ;
        RECT 194.200 75.200 194.500 111.800 ;
        RECT 195.000 85.800 195.400 86.200 ;
        RECT 194.200 74.800 194.600 75.200 ;
        RECT 193.400 72.800 193.800 73.200 ;
        RECT 195.000 66.200 195.300 85.800 ;
        RECT 195.000 65.800 195.400 66.200 ;
        RECT 192.600 49.800 193.000 50.200 ;
        RECT 195.800 46.200 196.100 133.800 ;
        RECT 196.600 129.800 197.000 130.200 ;
        RECT 195.800 45.800 196.200 46.200 ;
        RECT 165.400 41.800 165.800 42.200 ;
        RECT 171.000 41.800 171.400 42.200 ;
        RECT 187.000 42.100 187.400 42.200 ;
        RECT 186.200 41.800 187.400 42.100 ;
        RECT 190.200 41.800 190.600 42.200 ;
        RECT 164.600 36.800 165.000 37.200 ;
        RECT 171.000 29.200 171.300 41.800 ;
        RECT 179.800 29.800 180.200 30.200 ;
        RECT 171.000 28.800 171.400 29.200 ;
        RECT 171.800 28.800 172.200 29.200 ;
        RECT 171.800 26.200 172.100 28.800 ;
        RECT 179.800 27.200 180.100 29.800 ;
        RECT 179.800 26.800 180.200 27.200 ;
        RECT 163.800 25.800 164.200 26.200 ;
        RECT 171.800 25.800 172.200 26.200 ;
        RECT 163.000 13.800 163.400 14.200 ;
        RECT 163.800 11.200 164.100 25.800 ;
        RECT 186.200 25.200 186.500 41.800 ;
        RECT 196.600 31.200 196.900 129.800 ;
        RECT 197.400 33.200 197.700 133.800 ;
        RECT 198.200 130.100 198.600 130.200 ;
        RECT 199.000 130.100 199.300 135.800 ;
        RECT 198.200 129.800 199.300 130.100 ;
        RECT 197.400 32.800 197.800 33.200 ;
        RECT 196.600 30.800 197.000 31.200 ;
        RECT 199.800 26.200 200.100 140.800 ;
        RECT 202.200 137.800 202.600 138.200 ;
        RECT 202.200 128.200 202.500 137.800 ;
        RECT 202.200 127.800 202.600 128.200 ;
        RECT 202.200 127.200 202.500 127.800 ;
        RECT 202.200 126.800 202.600 127.200 ;
        RECT 200.600 102.800 201.000 103.200 ;
        RECT 200.600 57.200 200.900 102.800 ;
        RECT 201.400 86.800 201.800 87.200 ;
        RECT 201.400 86.200 201.700 86.800 ;
        RECT 201.400 85.800 201.800 86.200 ;
        RECT 201.400 68.800 201.800 69.200 ;
        RECT 201.400 68.200 201.700 68.800 ;
        RECT 201.400 67.800 201.800 68.200 ;
        RECT 201.400 65.800 201.800 66.200 ;
        RECT 200.600 56.800 201.000 57.200 ;
        RECT 201.400 48.200 201.700 65.800 ;
        RECT 202.200 52.800 202.600 53.200 ;
        RECT 201.400 47.800 201.800 48.200 ;
        RECT 202.200 47.200 202.500 52.800 ;
        RECT 202.200 46.800 202.600 47.200 ;
        RECT 199.800 25.800 200.200 26.200 ;
        RECT 186.200 24.800 186.600 25.200 ;
        RECT 163.800 10.800 164.200 11.200 ;
        RECT 157.400 9.800 157.800 10.200 ;
        RECT 121.400 6.800 121.800 7.200 ;
        RECT 29.400 5.800 29.800 6.200 ;
      LAYER via4 ;
        RECT 59.000 126.800 59.400 127.200 ;
        RECT 50.200 75.800 50.600 76.200 ;
        RECT 38.200 35.800 38.600 36.200 ;
        RECT 40.600 34.800 41.000 35.200 ;
        RECT 63.800 53.800 64.200 54.200 ;
        RECT 71.800 75.800 72.200 76.200 ;
        RECT 74.200 73.800 74.600 74.200 ;
        RECT 83.800 127.800 84.200 128.200 ;
        RECT 78.200 73.800 78.600 74.200 ;
        RECT 77.400 25.800 77.800 26.200 ;
        RECT 82.200 27.800 82.600 28.200 ;
        RECT 93.400 106.800 93.800 107.200 ;
        RECT 99.800 86.800 100.200 87.200 ;
        RECT 94.200 27.800 94.600 28.200 ;
        RECT 118.200 113.800 118.600 114.200 ;
        RECT 109.400 36.800 109.800 37.200 ;
        RECT 144.600 85.800 145.000 86.200 ;
        RECT 144.600 73.800 145.000 74.200 ;
        RECT 155.000 73.800 155.400 74.200 ;
        RECT 124.600 25.800 125.000 26.200 ;
        RECT 169.400 126.800 169.800 127.200 ;
        RECT 179.800 133.800 180.200 134.200 ;
        RECT 191.800 85.800 192.200 86.200 ;
      LAYER metal5 ;
        RECT 122.200 135.100 122.600 135.200 ;
        RECT 136.600 135.100 137.000 135.200 ;
        RECT 122.200 134.800 137.000 135.100 ;
        RECT 179.800 134.100 180.200 134.200 ;
        RECT 195.800 134.100 196.200 134.200 ;
        RECT 179.800 133.800 196.200 134.100 ;
        RECT 81.400 132.100 81.800 132.200 ;
        RECT 99.000 132.100 99.400 132.200 ;
        RECT 81.400 131.800 99.400 132.100 ;
        RECT 135.800 130.100 136.200 130.200 ;
        RECT 151.800 130.100 152.200 130.200 ;
        RECT 176.600 130.100 177.000 130.200 ;
        RECT 135.800 129.800 177.000 130.100 ;
        RECT 43.800 129.100 44.200 129.200 ;
        RECT 49.400 129.100 49.800 129.200 ;
        RECT 43.800 128.800 49.800 129.100 ;
        RECT 66.200 129.100 66.600 129.200 ;
        RECT 155.000 129.100 155.400 129.200 ;
        RECT 66.200 128.800 155.400 129.100 ;
        RECT 83.800 128.100 84.200 128.200 ;
        RECT 86.200 128.100 86.600 128.200 ;
        RECT 83.800 127.800 86.600 128.100 ;
        RECT 89.400 128.100 89.800 128.200 ;
        RECT 109.400 128.100 109.800 128.200 ;
        RECT 89.400 127.800 109.800 128.100 ;
        RECT 59.000 127.100 59.400 127.200 ;
        RECT 158.200 127.100 158.600 127.200 ;
        RECT 59.000 126.800 158.600 127.100 ;
        RECT 169.400 127.100 169.800 127.200 ;
        RECT 202.200 127.100 202.600 127.200 ;
        RECT 169.400 126.800 202.600 127.100 ;
        RECT 47.000 126.100 47.400 126.200 ;
        RECT 106.200 126.100 106.600 126.200 ;
        RECT 47.000 125.800 106.600 126.100 ;
        RECT 118.200 114.100 118.600 114.200 ;
        RECT 130.200 114.100 130.600 114.200 ;
        RECT 118.200 113.800 130.600 114.100 ;
        RECT 169.400 108.100 169.800 108.200 ;
        RECT 172.600 108.100 173.000 108.200 ;
        RECT 169.400 107.800 173.000 108.100 ;
        RECT 43.000 106.800 43.400 107.200 ;
        RECT 93.400 107.100 93.800 107.200 ;
        RECT 166.200 107.100 166.600 107.200 ;
        RECT 93.400 106.800 166.600 107.100 ;
        RECT 31.800 106.100 32.200 106.200 ;
        RECT 43.000 106.100 43.300 106.800 ;
        RECT 31.800 105.800 43.300 106.100 ;
        RECT 68.600 101.100 69.000 101.200 ;
        RECT 104.600 101.100 105.000 101.200 ;
        RECT 68.600 100.800 105.000 101.100 ;
        RECT 47.800 95.100 48.200 95.200 ;
        RECT 75.800 95.100 76.200 95.200 ;
        RECT 47.800 94.800 76.200 95.100 ;
        RECT 59.000 94.100 59.400 94.200 ;
        RECT 93.400 94.100 93.800 94.200 ;
        RECT 59.000 93.800 93.800 94.100 ;
        RECT 63.800 93.100 64.200 93.200 ;
        RECT 153.400 93.100 153.800 93.200 ;
        RECT 63.800 92.800 153.800 93.100 ;
        RECT 99.800 87.100 100.200 87.200 ;
        RECT 105.400 87.100 105.800 87.200 ;
        RECT 99.800 86.800 105.800 87.100 ;
        RECT 139.000 87.100 139.400 87.200 ;
        RECT 175.800 87.100 176.200 87.200 ;
        RECT 139.000 86.800 176.200 87.100 ;
        RECT 201.400 86.800 201.800 87.200 ;
        RECT 144.600 86.100 145.000 86.200 ;
        RECT 159.800 86.100 160.200 86.200 ;
        RECT 144.600 85.800 160.200 86.100 ;
        RECT 166.200 85.800 166.600 86.200 ;
        RECT 191.800 86.100 192.200 86.200 ;
        RECT 201.400 86.100 201.700 86.800 ;
        RECT 191.800 85.800 201.700 86.100 ;
        RECT 78.200 85.100 78.600 85.200 ;
        RECT 166.200 85.100 166.500 85.800 ;
        RECT 78.200 84.800 166.500 85.100 ;
        RECT 50.200 76.100 50.600 76.200 ;
        RECT 71.800 76.100 72.200 76.200 ;
        RECT 50.200 75.800 72.200 76.100 ;
        RECT 71.800 75.100 72.200 75.200 ;
        RECT 75.000 75.100 75.400 75.200 ;
        RECT 71.800 74.800 75.400 75.100 ;
        RECT 76.600 75.100 77.000 75.200 ;
        RECT 87.800 75.100 88.200 75.200 ;
        RECT 76.600 74.800 88.200 75.100 ;
        RECT 74.200 74.100 74.600 74.200 ;
        RECT 78.200 74.100 78.600 74.200 ;
        RECT 74.200 73.800 78.600 74.100 ;
        RECT 82.200 74.100 82.600 74.200 ;
        RECT 106.200 74.100 106.600 74.200 ;
        RECT 82.200 73.800 106.600 74.100 ;
        RECT 142.200 74.100 142.600 74.200 ;
        RECT 144.600 74.100 145.000 74.200 ;
        RECT 142.200 73.800 145.000 74.100 ;
        RECT 155.000 74.100 155.400 74.200 ;
        RECT 158.200 74.100 158.600 74.200 ;
        RECT 155.000 73.800 158.600 74.100 ;
        RECT 56.600 73.100 57.000 73.200 ;
        RECT 77.400 73.100 77.800 73.200 ;
        RECT 56.600 72.800 77.800 73.100 ;
        RECT 91.000 73.100 91.400 73.200 ;
        RECT 143.800 73.100 144.200 73.200 ;
        RECT 91.000 72.800 144.200 73.100 ;
        RECT 77.400 72.100 77.800 72.200 ;
        RECT 90.200 72.100 90.600 72.200 ;
        RECT 77.400 71.800 90.600 72.100 ;
        RECT 99.800 69.100 100.200 69.200 ;
        RECT 201.400 69.100 201.800 69.200 ;
        RECT 99.800 68.800 201.800 69.100 ;
        RECT 128.600 68.100 129.000 68.200 ;
        RECT 134.200 68.100 134.600 68.200 ;
        RECT 128.600 67.800 134.600 68.100 ;
        RECT 146.200 68.100 146.600 68.200 ;
        RECT 166.200 68.100 166.600 68.200 ;
        RECT 146.200 67.800 166.600 68.100 ;
        RECT 18.200 67.100 18.600 67.200 ;
        RECT 63.000 67.100 63.400 67.200 ;
        RECT 18.200 66.800 63.400 67.100 ;
        RECT 84.600 67.100 85.000 67.200 ;
        RECT 167.800 67.100 168.200 67.200 ;
        RECT 84.600 66.800 168.200 67.100 ;
        RECT 92.600 66.100 93.000 66.200 ;
        RECT 135.800 66.100 136.200 66.200 ;
        RECT 92.600 65.800 136.200 66.100 ;
        RECT 63.800 54.100 64.200 54.200 ;
        RECT 120.600 54.100 121.000 54.200 ;
        RECT 63.800 53.800 121.000 54.100 ;
        RECT 87.000 52.100 87.400 52.200 ;
        RECT 115.000 52.100 115.400 52.200 ;
        RECT 87.000 51.800 115.400 52.100 ;
        RECT 107.800 50.100 108.200 50.200 ;
        RECT 109.400 50.100 109.800 50.200 ;
        RECT 107.800 49.800 109.800 50.100 ;
        RECT 91.000 49.100 91.400 49.200 ;
        RECT 113.400 49.100 113.800 49.200 ;
        RECT 91.000 48.800 113.800 49.100 ;
        RECT 148.600 48.800 149.000 49.200 ;
        RECT 108.600 48.100 109.000 48.200 ;
        RECT 148.600 48.100 148.900 48.800 ;
        RECT 108.600 47.800 148.900 48.100 ;
        RECT 97.400 47.100 97.800 47.200 ;
        RECT 104.600 47.100 105.000 47.200 ;
        RECT 97.400 46.800 105.000 47.100 ;
        RECT 88.600 46.100 89.000 46.200 ;
        RECT 104.600 46.100 105.000 46.200 ;
        RECT 88.600 45.800 105.000 46.100 ;
        RECT 56.600 44.100 57.000 44.200 ;
        RECT 156.600 44.100 157.000 44.200 ;
        RECT 56.600 43.800 157.000 44.100 ;
        RECT 15.800 37.100 16.200 37.200 ;
        RECT 21.400 37.100 21.800 37.200 ;
        RECT 81.400 37.100 81.800 37.200 ;
        RECT 15.800 36.800 81.800 37.100 ;
        RECT 109.400 37.100 109.800 37.200 ;
        RECT 112.600 37.100 113.000 37.200 ;
        RECT 109.400 36.800 113.000 37.100 ;
        RECT 38.200 36.100 38.600 36.200 ;
        RECT 61.400 36.100 61.800 36.200 ;
        RECT 38.200 35.800 61.800 36.100 ;
        RECT 29.400 35.100 29.800 35.200 ;
        RECT 40.600 35.100 41.000 35.200 ;
        RECT 29.400 34.800 41.000 35.100 ;
        RECT 48.600 34.100 49.000 34.200 ;
        RECT 95.800 34.100 96.200 34.200 ;
        RECT 48.600 33.800 96.200 34.100 ;
        RECT 105.400 34.100 105.800 34.200 ;
        RECT 116.600 34.100 117.000 34.200 ;
        RECT 105.400 33.800 117.000 34.100 ;
        RECT 70.200 30.100 70.600 30.200 ;
        RECT 100.600 30.100 101.000 30.200 ;
        RECT 70.200 29.800 101.000 30.100 ;
        RECT 104.600 28.800 105.000 29.200 ;
        RECT 82.200 28.100 82.600 28.200 ;
        RECT 91.800 28.100 92.200 28.200 ;
        RECT 82.200 27.800 92.200 28.100 ;
        RECT 94.200 28.100 94.600 28.200 ;
        RECT 104.600 28.100 104.900 28.800 ;
        RECT 94.200 27.800 104.900 28.100 ;
        RECT 72.600 27.100 73.000 27.200 ;
        RECT 117.400 27.100 117.800 27.200 ;
        RECT 72.600 26.800 117.800 27.100 ;
        RECT 17.400 26.100 17.800 26.200 ;
        RECT 55.000 26.100 55.400 26.200 ;
        RECT 17.400 25.800 55.400 26.100 ;
        RECT 77.400 26.100 77.800 26.200 ;
        RECT 92.600 26.100 93.000 26.200 ;
        RECT 77.400 25.800 93.000 26.100 ;
        RECT 124.600 26.100 125.000 26.200 ;
        RECT 171.800 26.100 172.200 26.200 ;
        RECT 124.600 25.800 172.200 26.100 ;
        RECT 50.200 25.100 50.600 25.200 ;
        RECT 60.600 25.100 61.000 25.200 ;
        RECT 50.200 24.800 61.000 25.100 ;
  END
END fifo
END LIBRARY

