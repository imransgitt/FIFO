magic
tech scmos
timestamp 1713260442
<< metal1 >>
rect 496 1803 498 1807
rect 502 1803 505 1807
rect 509 1803 512 1807
rect 1528 1803 1530 1807
rect 1534 1803 1537 1807
rect 1541 1803 1544 1807
rect 1998 1768 2009 1771
rect 2006 1762 2009 1768
rect 190 1748 209 1751
rect 422 1748 457 1751
rect 1238 1748 1265 1751
rect 1974 1748 1985 1751
rect 2014 1748 2025 1751
rect 374 1741 377 1748
rect 374 1738 385 1741
rect 661 1738 662 1742
rect 850 1738 857 1741
rect 1142 1741 1145 1748
rect 1134 1738 1145 1741
rect 1298 1738 1313 1741
rect 2038 1738 2046 1741
rect 1086 1728 1094 1731
rect 1278 1728 1289 1731
rect 1016 1703 1018 1707
rect 1022 1703 1025 1707
rect 1029 1703 1032 1707
rect 662 1678 681 1681
rect 1118 1678 1134 1681
rect 538 1668 561 1671
rect 814 1668 822 1671
rect 1346 1668 1361 1671
rect 230 1658 233 1668
rect 606 1658 625 1661
rect 794 1658 801 1661
rect 814 1658 833 1661
rect 994 1658 1033 1661
rect 1074 1658 1081 1661
rect 1098 1658 1105 1661
rect 1110 1658 1118 1661
rect 1198 1658 1214 1661
rect 1230 1658 1238 1661
rect 1278 1658 1286 1661
rect 1838 1658 1857 1661
rect 1990 1658 1998 1661
rect 606 1648 609 1658
rect 814 1648 817 1658
rect 1854 1648 1857 1658
rect 842 1638 849 1641
rect 866 1638 869 1642
rect 1618 1638 1620 1642
rect 1998 1638 2017 1641
rect 2014 1628 2017 1638
rect 496 1603 498 1607
rect 502 1603 505 1607
rect 509 1603 512 1607
rect 1528 1603 1530 1607
rect 1534 1603 1537 1607
rect 1541 1603 1544 1607
rect 1797 1588 1798 1592
rect 973 1568 974 1572
rect 530 1558 534 1562
rect 542 1558 561 1561
rect 86 1548 102 1551
rect 522 1548 529 1551
rect 598 1542 601 1551
rect 726 1551 729 1561
rect 942 1558 958 1561
rect 1238 1558 1246 1561
rect 1850 1558 1854 1562
rect 1862 1558 1870 1561
rect 726 1548 745 1551
rect 974 1548 990 1551
rect 1582 1548 1585 1558
rect 1798 1548 1817 1551
rect 1054 1538 1070 1541
rect 1150 1538 1153 1548
rect 142 1531 146 1533
rect 142 1528 150 1531
rect 374 1528 393 1531
rect 1010 1528 1033 1531
rect 1082 1528 1097 1531
rect 1162 1528 1177 1531
rect 1016 1503 1018 1507
rect 1022 1503 1025 1507
rect 1029 1503 1032 1507
rect 1898 1488 1899 1492
rect 1970 1488 1972 1492
rect 662 1478 670 1481
rect 1110 1478 1126 1481
rect 1956 1478 1958 1482
rect 398 1472 402 1474
rect 138 1468 145 1471
rect 174 1468 182 1471
rect 918 1471 922 1474
rect 910 1468 922 1471
rect 1006 1468 1014 1471
rect 350 1458 366 1461
rect 446 1458 462 1461
rect 550 1458 569 1461
rect 886 1458 905 1461
rect 962 1458 977 1461
rect 1430 1461 1433 1471
rect 1614 1468 1625 1471
rect 1702 1468 1710 1471
rect 1738 1468 1753 1471
rect 1758 1468 1774 1471
rect 1806 1468 1822 1471
rect 1430 1458 1449 1461
rect 1478 1458 1486 1461
rect 1510 1458 1537 1461
rect 1566 1458 1585 1461
rect 1630 1458 1657 1461
rect 1662 1458 1681 1461
rect 1890 1458 1897 1461
rect 1902 1458 1921 1461
rect 566 1448 569 1458
rect 886 1448 889 1458
rect 1054 1456 1058 1458
rect 1270 1456 1274 1458
rect 1054 1448 1062 1451
rect 1174 1442 1177 1451
rect 1466 1448 1473 1451
rect 1478 1448 1481 1458
rect 1902 1448 1905 1458
rect 1805 1438 1806 1442
rect 1926 1438 1950 1441
rect 1070 1428 1073 1438
rect 502 1418 518 1421
rect 1314 1418 1315 1422
rect 496 1403 498 1407
rect 502 1403 505 1407
rect 509 1403 512 1407
rect 1528 1403 1530 1407
rect 1534 1403 1537 1407
rect 1541 1403 1544 1407
rect 614 1368 622 1371
rect 646 1351 649 1361
rect 630 1348 649 1351
rect 674 1348 689 1351
rect 790 1351 793 1361
rect 774 1348 793 1351
rect 942 1351 945 1361
rect 926 1348 945 1351
rect 998 1348 1022 1351
rect 1126 1351 1129 1361
rect 1806 1358 1817 1361
rect 1806 1352 1809 1358
rect 1126 1348 1145 1351
rect 1306 1348 1313 1351
rect 1462 1348 1473 1351
rect 1550 1348 1566 1351
rect 1642 1348 1649 1351
rect 1722 1348 1737 1351
rect 1794 1348 1801 1351
rect 1462 1342 1465 1348
rect 494 1338 518 1341
rect 1038 1338 1046 1341
rect 1274 1338 1281 1341
rect 1798 1338 1806 1341
rect 1870 1338 1889 1341
rect 1962 1338 1969 1341
rect 2038 1338 2046 1341
rect 1290 1328 1305 1331
rect 1342 1331 1345 1338
rect 1334 1328 1345 1331
rect 1606 1331 1610 1333
rect 1358 1328 1377 1331
rect 1606 1328 1614 1331
rect 717 1318 718 1322
rect 1074 1318 1075 1322
rect 1016 1303 1018 1307
rect 1022 1303 1025 1307
rect 1029 1303 1032 1307
rect 426 1288 427 1292
rect 94 1278 105 1281
rect 594 1278 598 1282
rect 886 1278 898 1281
rect 94 1277 98 1278
rect 894 1277 898 1278
rect 310 1262 313 1271
rect 1010 1268 1033 1271
rect 1126 1268 1145 1271
rect 1270 1268 1282 1271
rect 1430 1271 1433 1281
rect 1546 1278 1561 1281
rect 1566 1278 1585 1281
rect 1702 1278 1713 1281
rect 1426 1268 1433 1271
rect 1586 1268 1593 1271
rect 1618 1268 1625 1271
rect 38 1258 54 1261
rect 286 1258 305 1261
rect 350 1258 358 1261
rect 522 1258 529 1261
rect 778 1258 785 1261
rect 998 1258 1033 1261
rect 1398 1258 1417 1261
rect 1670 1262 1673 1271
rect 1862 1268 1870 1271
rect 1958 1268 1974 1271
rect 1674 1258 1681 1261
rect 1922 1258 1929 1261
rect 1962 1258 1977 1261
rect 2038 1258 2046 1261
rect 274 1248 278 1252
rect 286 1248 289 1258
rect 570 1248 574 1252
rect 1030 1248 1033 1258
rect 1398 1248 1401 1258
rect 406 1238 414 1241
rect 1202 1238 1205 1242
rect 1347 1238 1350 1242
rect 1170 1228 1171 1232
rect 837 1218 838 1222
rect 861 1218 862 1222
rect 496 1203 498 1207
rect 502 1203 505 1207
rect 509 1203 512 1207
rect 1528 1203 1530 1207
rect 1534 1203 1537 1207
rect 1541 1203 1544 1207
rect 1146 1188 1148 1192
rect 1229 1188 1230 1192
rect 1658 1188 1659 1192
rect 1293 1178 1294 1182
rect 171 1168 174 1172
rect 350 1168 358 1171
rect 38 1148 54 1151
rect 134 1148 142 1151
rect 202 1148 209 1151
rect 382 1151 385 1161
rect 366 1148 385 1151
rect 502 1148 510 1151
rect 514 1148 526 1151
rect 550 1151 553 1161
rect 894 1158 913 1161
rect 550 1148 569 1151
rect 606 1148 614 1151
rect 766 1148 774 1151
rect 798 1148 809 1151
rect 862 1148 870 1151
rect 958 1148 966 1151
rect 1062 1151 1065 1161
rect 1270 1158 1281 1161
rect 1046 1148 1065 1151
rect 1230 1148 1238 1151
rect 798 1142 801 1148
rect 482 1138 489 1141
rect 574 1138 582 1141
rect 746 1138 753 1141
rect 834 1138 849 1141
rect 866 1138 873 1141
rect 1026 1138 1041 1141
rect 1110 1138 1118 1141
rect 1318 1138 1326 1141
rect 1942 1138 1954 1141
rect 190 1131 194 1133
rect 190 1128 201 1131
rect 438 1128 449 1131
rect 1546 1128 1553 1131
rect 1014 1118 1022 1121
rect 1016 1103 1018 1107
rect 1022 1103 1025 1107
rect 1029 1103 1032 1107
rect 1270 1078 1281 1081
rect 1286 1078 1305 1081
rect 1390 1078 1402 1081
rect 1270 1077 1274 1078
rect 1398 1077 1402 1078
rect 1630 1078 1649 1081
rect 1766 1078 1778 1081
rect 1598 1077 1602 1078
rect 166 1068 174 1071
rect 466 1068 473 1071
rect 618 1068 625 1071
rect 894 1068 905 1071
rect 1366 1068 1374 1071
rect 1486 1068 1514 1071
rect 1654 1071 1657 1078
rect 1774 1077 1778 1078
rect 1654 1068 1673 1071
rect 2038 1068 2046 1071
rect 142 1058 161 1061
rect 170 1058 174 1061
rect 178 1058 185 1061
rect 230 1058 249 1061
rect 254 1058 262 1061
rect 322 1058 329 1061
rect 370 1058 377 1061
rect 486 1058 510 1061
rect 790 1058 798 1061
rect 854 1061 857 1068
rect 894 1062 897 1068
rect 854 1058 865 1061
rect 990 1058 1025 1061
rect 1542 1058 1558 1061
rect 1742 1058 1761 1061
rect 1950 1058 1958 1061
rect 1970 1058 1977 1061
rect 1990 1058 2009 1061
rect 130 1048 134 1052
rect 142 1048 145 1058
rect 310 1048 321 1051
rect 390 1048 401 1051
rect 1022 1048 1025 1058
rect 1990 1048 1993 1058
rect 746 1018 747 1022
rect 885 1018 886 1022
rect 496 1003 498 1007
rect 502 1003 505 1007
rect 509 1003 512 1007
rect 1528 1003 1530 1007
rect 1534 1003 1537 1007
rect 1541 1003 1544 1007
rect 813 978 814 982
rect 1722 968 1723 972
rect 1858 968 1861 972
rect 198 958 217 961
rect 570 958 574 962
rect 110 948 118 951
rect 226 948 233 951
rect 334 948 342 951
rect 378 948 385 951
rect 550 948 558 951
rect 586 948 593 951
rect 762 948 777 951
rect 814 948 830 951
rect 950 948 958 951
rect 1198 951 1201 961
rect 1182 948 1201 951
rect 1214 948 1222 951
rect 1646 951 1649 961
rect 1734 958 1745 961
rect 1630 948 1649 951
rect 282 938 289 941
rect 502 938 510 941
rect 606 938 625 941
rect 894 938 902 941
rect 958 938 966 941
rect 1002 938 1009 941
rect 1194 938 1201 941
rect 1494 938 1502 941
rect 1582 938 1601 941
rect 1618 938 1625 941
rect 166 936 170 938
rect 398 928 409 931
rect 622 928 625 938
rect 1414 928 1433 931
rect 1438 928 1441 938
rect 1546 928 1561 931
rect 1582 928 1585 938
rect 1838 931 1842 933
rect 1950 931 1954 933
rect 1830 928 1842 931
rect 1942 928 1954 931
rect 1016 903 1018 907
rect 1022 903 1025 907
rect 1029 903 1032 907
rect 334 878 345 881
rect 350 878 369 881
rect 470 878 498 881
rect 1294 878 1313 881
rect 1606 878 1618 881
rect 1950 878 1962 881
rect 334 877 338 878
rect 494 877 498 878
rect 1614 877 1618 878
rect 1958 877 1962 878
rect 1062 872 1066 874
rect 122 868 129 871
rect 150 868 158 871
rect 298 868 299 872
rect 610 868 617 871
rect 1101 868 1102 872
rect 1314 868 1321 871
rect 1326 868 1334 871
rect 1534 868 1566 871
rect 1594 868 1601 871
rect 1886 868 1894 871
rect 110 858 129 861
rect 342 861 345 868
rect 334 858 345 861
rect 446 858 465 861
rect 598 858 617 861
rect 674 858 681 861
rect 726 858 734 861
rect 810 858 817 861
rect 874 858 882 861
rect 958 858 977 861
rect 998 858 1033 861
rect 1106 858 1121 861
rect 1770 858 1777 861
rect 126 848 129 858
rect 334 857 338 858
rect 206 848 217 851
rect 422 848 433 851
rect 614 848 617 858
rect 678 848 681 858
rect 1030 848 1033 858
rect 1722 848 1726 852
rect 1750 848 1769 851
rect 725 828 726 832
rect 957 818 958 822
rect 1485 818 1486 822
rect 496 803 498 807
rect 502 803 505 807
rect 509 803 512 807
rect 1528 803 1530 807
rect 1534 803 1537 807
rect 1541 803 1544 807
rect 730 788 731 792
rect 1146 788 1147 792
rect 538 778 539 782
rect 414 768 422 771
rect 1834 768 1837 772
rect 38 748 46 751
rect 162 748 169 751
rect 174 748 182 751
rect 446 751 449 761
rect 506 758 513 761
rect 430 748 449 751
rect 550 751 553 758
rect 530 748 537 751
rect 550 748 561 751
rect 598 748 609 751
rect 638 748 654 751
rect 682 748 694 751
rect 842 748 849 751
rect 1102 751 1105 761
rect 1086 748 1105 751
rect 1190 751 1194 753
rect 1162 748 1169 751
rect 1174 748 1194 751
rect 94 731 98 733
rect 246 732 249 742
rect 442 738 449 741
rect 558 741 561 748
rect 606 742 609 748
rect 514 738 529 741
rect 558 738 569 741
rect 710 738 713 748
rect 1390 751 1393 761
rect 1390 748 1409 751
rect 1750 748 1758 751
rect 1866 748 1873 751
rect 2010 748 2017 751
rect 1786 738 1793 741
rect 982 733 986 738
rect 94 728 105 731
rect 110 728 129 731
rect 862 728 873 731
rect 950 728 958 731
rect 1286 728 1289 738
rect 1974 732 1978 736
rect 1318 728 1337 731
rect 1646 728 1665 731
rect 1766 728 1785 731
rect 298 718 299 722
rect 1016 703 1018 707
rect 1022 703 1025 707
rect 1029 703 1032 707
rect 694 677 698 678
rect 430 672 434 674
rect 138 668 145 671
rect 726 671 729 681
rect 1214 678 1230 681
rect 1710 678 1722 681
rect 1886 678 1897 681
rect 1214 674 1218 678
rect 1630 674 1634 678
rect 1718 677 1722 678
rect 726 668 745 671
rect 806 668 817 671
rect 894 668 905 671
rect 950 668 961 671
rect 1006 668 1030 671
rect 1198 671 1202 674
rect 1194 668 1202 671
rect 1430 668 1441 671
rect 1482 668 1489 671
rect 1694 668 1705 671
rect 1806 668 1814 671
rect 38 658 46 661
rect 118 658 134 661
rect 302 658 318 661
rect 514 658 529 661
rect 638 658 654 661
rect 830 658 846 661
rect 974 658 993 661
rect 1022 658 1049 661
rect 1318 658 1326 661
rect 1334 658 1353 661
rect 1438 661 1441 668
rect 1438 658 1446 661
rect 1694 662 1697 668
rect 1762 658 1777 661
rect 1922 658 1937 661
rect 1022 652 1025 658
rect 1350 648 1353 658
rect 1446 648 1449 658
rect 1534 648 1542 651
rect 326 638 334 641
rect 411 638 414 642
rect 530 638 531 642
rect 496 603 498 607
rect 502 603 505 607
rect 509 603 512 607
rect 1528 603 1530 607
rect 1534 603 1537 607
rect 1541 603 1544 607
rect 418 588 419 592
rect 621 588 622 592
rect 869 588 870 592
rect 1069 588 1070 592
rect 210 568 211 572
rect 342 568 350 571
rect 562 568 563 572
rect 134 548 142 551
rect 222 551 225 561
rect 202 548 209 551
rect 222 548 241 551
rect 286 548 294 551
rect 374 551 377 561
rect 358 548 377 551
rect 574 551 577 561
rect 778 558 782 562
rect 574 548 593 551
rect 634 548 641 551
rect 790 551 793 561
rect 790 548 809 551
rect 910 551 913 561
rect 1050 558 1057 561
rect 910 548 929 551
rect 1126 551 1129 561
rect 1070 548 1089 551
rect 1110 548 1129 551
rect 1242 548 1249 551
rect 1310 551 1313 561
rect 1310 548 1329 551
rect 1590 551 1593 558
rect 1582 548 1593 551
rect 1726 548 1734 551
rect 1938 548 1945 551
rect 1994 548 2009 551
rect 342 538 353 541
rect 538 538 550 541
rect 910 538 918 541
rect 1094 538 1102 541
rect 1558 538 1566 541
rect 1946 538 1953 541
rect 342 536 346 538
rect 1094 528 1097 538
rect 1414 533 1418 538
rect 1598 531 1602 533
rect 1590 528 1602 531
rect 1894 531 1898 533
rect 1766 528 1777 531
rect 1894 528 1905 531
rect 1966 528 1985 531
rect 1016 503 1018 507
rect 1022 503 1025 507
rect 1029 503 1032 507
rect 86 478 105 481
rect 458 478 474 481
rect 470 474 474 478
rect 790 478 801 481
rect 1178 478 1186 481
rect 1446 478 1465 481
rect 1638 478 1649 481
rect 1838 478 1849 481
rect 1882 478 1883 482
rect 790 477 794 478
rect 1182 477 1186 478
rect 1838 477 1842 478
rect 1990 472 1994 474
rect 118 468 126 471
rect 182 468 190 471
rect 214 468 222 471
rect 998 468 1006 471
rect 1122 468 1129 471
rect 142 458 161 461
rect 186 458 201 461
rect 214 458 233 461
rect 366 458 385 461
rect 1278 462 1281 471
rect 1306 468 1321 471
rect 1718 468 1726 471
rect 2026 468 2041 471
rect 450 458 457 461
rect 526 458 553 461
rect 638 458 654 461
rect 734 458 750 461
rect 1226 458 1241 461
rect 1462 458 1465 468
rect 1562 458 1569 461
rect 1662 458 1670 461
rect 1894 458 1902 461
rect 1942 458 1958 461
rect 158 448 161 458
rect 214 448 217 458
rect 366 448 369 458
rect 1694 448 1702 451
rect 1979 438 1982 442
rect 496 403 498 407
rect 502 403 505 407
rect 509 403 512 407
rect 1528 403 1530 407
rect 1534 403 1537 407
rect 1541 403 1544 407
rect 442 388 443 392
rect 554 388 555 392
rect 1366 368 1374 371
rect 1402 368 1405 372
rect 350 358 369 361
rect 10 348 17 351
rect 214 348 222 351
rect 262 348 270 351
rect 590 351 593 358
rect 582 348 593 351
rect 606 348 614 351
rect 678 351 681 361
rect 678 348 697 351
rect 862 351 865 361
rect 1782 358 1790 361
rect 862 348 881 351
rect 938 348 953 351
rect 1210 348 1225 351
rect 1310 348 1326 351
rect 1426 348 1441 351
rect 1626 348 1641 351
rect 1898 348 1913 351
rect 170 338 177 341
rect 582 338 593 341
rect 626 338 633 341
rect 886 338 898 341
rect 998 338 1033 341
rect 1150 338 1158 341
rect 1542 338 1550 341
rect 1766 338 1774 341
rect 1850 338 1858 341
rect 582 332 585 338
rect 894 336 898 338
rect 1854 336 1858 338
rect 1166 331 1170 333
rect 1158 328 1170 331
rect 1382 331 1386 333
rect 1582 331 1586 333
rect 1270 328 1289 331
rect 1374 328 1386 331
rect 1574 328 1586 331
rect 1686 328 1705 331
rect 1806 328 1825 331
rect 1016 303 1018 307
rect 1022 303 1025 307
rect 1029 303 1032 307
rect 574 278 585 281
rect 622 278 633 281
rect 190 268 202 271
rect 286 271 290 274
rect 630 272 633 278
rect 286 268 297 271
rect 506 268 529 271
rect 1078 271 1081 281
rect 1086 278 1105 281
rect 1286 278 1297 281
rect 1326 272 1330 274
rect 1066 268 1081 271
rect 1130 268 1137 271
rect 1226 268 1233 271
rect 1582 271 1585 281
rect 1790 274 1794 278
rect 1582 268 1601 271
rect 302 258 321 261
rect 470 258 489 261
rect 654 258 662 261
rect 718 258 726 261
rect 790 258 809 261
rect 834 258 849 261
rect 966 258 974 261
rect 1182 258 1190 261
rect 1202 258 1209 261
rect 1370 258 1385 261
rect 1478 258 1486 261
rect 1546 258 1558 261
rect 1662 258 1670 261
rect 1722 258 1737 261
rect 1946 258 1953 261
rect 318 248 321 258
rect 458 248 462 252
rect 470 248 473 258
rect 650 248 654 252
rect 714 248 718 252
rect 806 248 809 258
rect 1466 238 1469 242
rect 1698 238 1701 242
rect 1181 218 1182 222
rect 1970 218 1971 222
rect 2038 218 2046 221
rect 496 203 498 207
rect 502 203 505 207
rect 509 203 512 207
rect 1528 203 1530 207
rect 1534 203 1537 207
rect 1541 203 1544 207
rect 1490 168 1493 172
rect 38 148 54 151
rect 210 148 217 151
rect 278 151 281 161
rect 278 148 297 151
rect 334 151 337 161
rect 334 148 353 151
rect 542 151 545 161
rect 542 148 561 151
rect 590 148 598 151
rect 606 148 617 151
rect 94 138 102 141
rect 382 138 385 148
rect 614 142 617 148
rect 806 148 814 151
rect 862 151 865 161
rect 846 148 865 151
rect 926 148 942 151
rect 998 148 1017 151
rect 1166 151 1169 161
rect 1150 148 1169 151
rect 998 142 1001 148
rect 1398 148 1414 151
rect 1514 148 1529 151
rect 2010 148 2017 151
rect 774 138 785 141
rect 94 136 98 138
rect 982 132 986 133
rect 126 128 145 131
rect 1270 131 1274 136
rect 1258 128 1274 131
rect 1422 128 1441 131
rect 1570 128 1585 131
rect 1590 128 1609 131
rect 1646 128 1665 131
rect 1774 128 1793 131
rect 1830 128 1849 131
rect 2030 118 2038 121
rect 1016 103 1018 107
rect 1022 103 1025 107
rect 1029 103 1032 107
rect 238 78 246 81
rect 254 78 273 81
rect 238 77 242 78
rect 518 68 546 71
rect 598 68 601 78
rect 614 74 618 78
rect 630 71 634 74
rect 822 72 826 74
rect 630 68 641 71
rect 658 68 665 71
rect 1138 68 1145 71
rect 1198 71 1201 81
rect 1334 78 1346 81
rect 1342 77 1346 78
rect 1182 68 1201 71
rect 1374 68 1377 78
rect 2006 72 2010 74
rect 1918 68 1930 71
rect 270 58 273 68
rect 646 58 665 61
rect 726 58 742 61
rect 1126 58 1145 61
rect 1274 58 1289 61
rect 1394 58 1401 61
rect 1682 58 1697 61
rect 1874 58 1889 61
rect 410 48 414 52
rect 662 48 665 58
rect 1142 48 1145 58
rect 496 3 498 7
rect 502 3 505 7
rect 509 3 512 7
rect 1528 3 1530 7
rect 1534 3 1537 7
rect 1541 3 1544 7
<< m2contact >>
rect 498 1803 502 1807
rect 505 1803 509 1807
rect 1530 1803 1534 1807
rect 1537 1803 1541 1807
rect 6 1788 10 1792
rect 30 1788 34 1792
rect 174 1788 178 1792
rect 350 1788 354 1792
rect 598 1788 602 1792
rect 1454 1788 1458 1792
rect 1510 1788 1514 1792
rect 1758 1788 1762 1792
rect 958 1779 962 1783
rect 1950 1768 1954 1772
rect 350 1758 354 1762
rect 598 1758 602 1762
rect 958 1756 962 1760
rect 1454 1758 1458 1762
rect 1510 1758 1514 1762
rect 1758 1758 1762 1762
rect 1934 1758 1938 1762
rect 2006 1758 2010 1762
rect 22 1748 26 1752
rect 46 1748 50 1752
rect 142 1748 146 1752
rect 166 1748 170 1752
rect 334 1748 338 1752
rect 350 1748 354 1752
rect 374 1748 378 1752
rect 398 1748 402 1752
rect 494 1748 498 1752
rect 678 1748 682 1752
rect 774 1748 778 1752
rect 942 1748 946 1752
rect 1118 1748 1122 1752
rect 1142 1748 1146 1752
rect 1350 1748 1354 1752
rect 1462 1748 1466 1752
rect 1510 1748 1514 1752
rect 1614 1748 1618 1752
rect 1774 1748 1778 1752
rect 1942 1748 1946 1752
rect 54 1738 58 1742
rect 126 1738 130 1742
rect 150 1738 154 1742
rect 302 1738 306 1742
rect 550 1738 554 1742
rect 662 1738 666 1742
rect 702 1738 706 1742
rect 750 1738 754 1742
rect 798 1738 802 1742
rect 814 1738 818 1742
rect 846 1738 850 1742
rect 918 1738 922 1742
rect 990 1738 994 1742
rect 1150 1738 1154 1742
rect 1214 1738 1218 1742
rect 1294 1738 1298 1742
rect 1406 1738 1410 1742
rect 1558 1738 1562 1742
rect 1670 1738 1674 1742
rect 1734 1738 1738 1742
rect 1806 1738 1810 1742
rect 2046 1738 2050 1742
rect 286 1728 290 1732
rect 534 1728 538 1732
rect 1006 1728 1010 1732
rect 1094 1728 1098 1732
rect 1222 1728 1226 1732
rect 1254 1728 1258 1732
rect 1390 1728 1394 1732
rect 1574 1728 1578 1732
rect 1822 1728 1826 1732
rect 1926 1728 1930 1732
rect 1950 1728 1954 1732
rect 1966 1728 1970 1732
rect 2006 1728 2010 1732
rect 110 1718 114 1722
rect 406 1718 410 1722
rect 622 1718 626 1722
rect 718 1718 722 1722
rect 822 1718 826 1722
rect 1230 1718 1234 1722
rect 1270 1718 1274 1722
rect 1286 1718 1290 1722
rect 1654 1718 1658 1722
rect 1902 1718 1906 1722
rect 1918 1718 1922 1722
rect 1018 1703 1022 1707
rect 1025 1703 1029 1707
rect 14 1688 18 1692
rect 190 1688 194 1692
rect 366 1688 370 1692
rect 606 1688 610 1692
rect 654 1688 658 1692
rect 966 1688 970 1692
rect 1262 1688 1266 1692
rect 1566 1688 1570 1692
rect 1854 1688 1858 1692
rect 1942 1688 1946 1692
rect 94 1678 98 1682
rect 270 1678 274 1682
rect 446 1678 450 1682
rect 686 1678 690 1682
rect 1046 1678 1050 1682
rect 1094 1678 1098 1682
rect 1214 1678 1218 1682
rect 1238 1678 1242 1682
rect 1438 1678 1442 1682
rect 1734 1678 1738 1682
rect 1902 1678 1906 1682
rect 1910 1678 1914 1682
rect 2038 1678 2042 1682
rect 2046 1678 2050 1682
rect 110 1668 114 1672
rect 230 1668 234 1672
rect 286 1668 290 1672
rect 462 1668 466 1672
rect 534 1668 538 1672
rect 582 1668 586 1672
rect 630 1668 634 1672
rect 646 1668 650 1672
rect 702 1668 706 1672
rect 790 1668 794 1672
rect 822 1668 826 1672
rect 838 1668 842 1672
rect 926 1668 930 1672
rect 942 1668 946 1672
rect 990 1668 994 1672
rect 1006 1668 1010 1672
rect 1054 1668 1058 1672
rect 1142 1668 1146 1672
rect 1182 1668 1186 1672
rect 1286 1668 1290 1672
rect 1294 1668 1298 1672
rect 1342 1668 1346 1672
rect 1454 1668 1458 1672
rect 1542 1668 1546 1672
rect 1590 1668 1594 1672
rect 1598 1668 1602 1672
rect 1646 1668 1650 1672
rect 1718 1668 1722 1672
rect 1830 1668 1834 1672
rect 1878 1668 1882 1672
rect 1894 1668 1898 1672
rect 1918 1668 1922 1672
rect 1966 1668 1970 1672
rect 1974 1668 1978 1672
rect 158 1658 162 1662
rect 334 1658 338 1662
rect 510 1658 514 1662
rect 574 1658 578 1662
rect 590 1658 594 1662
rect 638 1658 642 1662
rect 670 1658 674 1662
rect 718 1659 722 1663
rect 750 1658 754 1662
rect 790 1658 794 1662
rect 902 1658 906 1662
rect 990 1658 994 1662
rect 1070 1658 1074 1662
rect 1094 1658 1098 1662
rect 1118 1658 1122 1662
rect 1158 1658 1162 1662
rect 1190 1658 1194 1662
rect 1214 1658 1218 1662
rect 1238 1658 1242 1662
rect 1254 1658 1258 1662
rect 1286 1658 1290 1662
rect 1486 1658 1490 1662
rect 1670 1658 1674 1662
rect 1774 1658 1778 1662
rect 1870 1658 1874 1662
rect 1886 1658 1890 1662
rect 1982 1658 1986 1662
rect 1998 1658 2002 1662
rect 2014 1658 2018 1662
rect 158 1648 162 1652
rect 318 1650 322 1654
rect 494 1650 498 1654
rect 614 1648 618 1652
rect 822 1648 826 1652
rect 1062 1648 1066 1652
rect 1070 1648 1074 1652
rect 1086 1648 1090 1652
rect 1126 1648 1130 1652
rect 1150 1648 1154 1652
rect 1206 1648 1210 1652
rect 1246 1648 1250 1652
rect 1262 1648 1266 1652
rect 1502 1648 1506 1652
rect 1670 1648 1674 1652
rect 1846 1648 1850 1652
rect 2006 1648 2010 1652
rect 838 1638 842 1642
rect 862 1638 866 1642
rect 1166 1638 1170 1642
rect 1318 1638 1322 1642
rect 1614 1638 1618 1642
rect 2022 1638 2026 1642
rect 494 1627 498 1631
rect 158 1618 162 1622
rect 318 1618 322 1622
rect 558 1618 562 1622
rect 782 1618 786 1622
rect 1030 1618 1034 1622
rect 1158 1618 1162 1622
rect 1230 1618 1234 1622
rect 1502 1618 1506 1622
rect 1670 1618 1674 1622
rect 1814 1618 1818 1622
rect 498 1603 502 1607
rect 505 1603 509 1607
rect 1530 1603 1534 1607
rect 1537 1603 1541 1607
rect 326 1588 330 1592
rect 798 1588 802 1592
rect 1038 1588 1042 1592
rect 1398 1588 1402 1592
rect 1574 1588 1578 1592
rect 1630 1588 1634 1592
rect 1798 1588 1802 1592
rect 6 1568 10 1572
rect 30 1568 34 1572
rect 974 1568 978 1572
rect 326 1558 330 1562
rect 526 1558 530 1562
rect 566 1558 570 1562
rect 22 1548 26 1552
rect 46 1548 50 1552
rect 102 1548 106 1552
rect 166 1548 170 1552
rect 181 1548 185 1552
rect 334 1548 338 1552
rect 350 1548 354 1552
rect 382 1548 386 1552
rect 438 1548 442 1552
rect 518 1548 522 1552
rect 574 1548 578 1552
rect 630 1547 634 1551
rect 662 1548 666 1552
rect 710 1548 714 1552
rect 718 1548 722 1552
rect 734 1558 738 1562
rect 774 1558 778 1562
rect 798 1558 802 1562
rect 958 1558 962 1562
rect 1086 1558 1090 1562
rect 1166 1558 1170 1562
rect 1214 1558 1218 1562
rect 1246 1558 1250 1562
rect 1398 1558 1402 1562
rect 1574 1558 1578 1562
rect 1582 1558 1586 1562
rect 1630 1558 1634 1562
rect 1846 1558 1850 1562
rect 1870 1558 1874 1562
rect 1910 1558 1914 1562
rect 814 1548 818 1552
rect 902 1548 906 1552
rect 990 1548 994 1552
rect 1062 1548 1066 1552
rect 1110 1548 1114 1552
rect 1118 1548 1122 1552
rect 1150 1548 1154 1552
rect 1190 1548 1194 1552
rect 1382 1548 1386 1552
rect 1470 1548 1474 1552
rect 1630 1548 1634 1552
rect 1790 1548 1794 1552
rect 1846 1548 1850 1552
rect 1894 1548 1898 1552
rect 1902 1548 1906 1552
rect 1934 1548 1938 1552
rect 1982 1548 1986 1552
rect 62 1538 66 1542
rect 94 1538 98 1542
rect 278 1538 282 1542
rect 358 1538 362 1542
rect 446 1538 450 1542
rect 518 1538 522 1542
rect 550 1538 554 1542
rect 582 1538 586 1542
rect 598 1538 602 1542
rect 702 1538 706 1542
rect 750 1538 754 1542
rect 758 1538 762 1542
rect 766 1538 770 1542
rect 846 1538 850 1542
rect 982 1538 986 1542
rect 1070 1538 1074 1542
rect 1198 1538 1202 1542
rect 1222 1538 1226 1542
rect 1350 1538 1354 1542
rect 1526 1538 1530 1542
rect 1678 1538 1682 1542
rect 1838 1538 1842 1542
rect 1886 1538 1890 1542
rect 1942 1538 1946 1542
rect 1958 1538 1962 1542
rect 150 1528 154 1532
rect 262 1528 266 1532
rect 398 1528 402 1532
rect 598 1528 602 1532
rect 862 1528 866 1532
rect 1006 1528 1010 1532
rect 1046 1528 1050 1532
rect 1102 1528 1106 1532
rect 1134 1528 1138 1532
rect 1334 1528 1338 1532
rect 1510 1528 1514 1532
rect 1694 1528 1698 1532
rect 1806 1528 1810 1532
rect 1830 1528 1834 1532
rect 1870 1528 1874 1532
rect 158 1518 162 1522
rect 366 1518 370 1522
rect 494 1518 498 1522
rect 694 1518 698 1522
rect 998 1518 1002 1522
rect 1182 1518 1186 1522
rect 1214 1518 1218 1522
rect 1238 1518 1242 1522
rect 1254 1518 1258 1522
rect 1430 1518 1434 1522
rect 1774 1518 1778 1522
rect 1822 1518 1826 1522
rect 1878 1518 1882 1522
rect 1918 1518 1922 1522
rect 2038 1518 2042 1522
rect 1018 1503 1022 1507
rect 1025 1503 1029 1507
rect 94 1488 98 1492
rect 150 1488 154 1492
rect 614 1488 618 1492
rect 654 1488 658 1492
rect 1334 1488 1338 1492
rect 1406 1488 1410 1492
rect 1550 1488 1554 1492
rect 1694 1488 1698 1492
rect 1838 1488 1842 1492
rect 1894 1488 1898 1492
rect 1966 1488 1970 1492
rect 1998 1488 2002 1492
rect 158 1478 162 1482
rect 534 1478 538 1482
rect 630 1478 634 1482
rect 670 1478 674 1482
rect 758 1478 762 1482
rect 846 1478 850 1482
rect 1302 1478 1306 1482
rect 1358 1478 1362 1482
rect 1510 1478 1514 1482
rect 1606 1478 1610 1482
rect 1742 1478 1746 1482
rect 1814 1478 1818 1482
rect 1878 1478 1882 1482
rect 1910 1478 1914 1482
rect 1958 1478 1962 1482
rect 30 1468 34 1472
rect 102 1468 106 1472
rect 118 1468 122 1472
rect 134 1468 138 1472
rect 166 1468 170 1472
rect 182 1468 186 1472
rect 198 1468 202 1472
rect 214 1468 218 1472
rect 230 1468 234 1472
rect 358 1468 362 1472
rect 398 1468 402 1472
rect 446 1468 450 1472
rect 542 1468 546 1472
rect 566 1468 570 1472
rect 590 1468 594 1472
rect 774 1468 778 1472
rect 862 1468 866 1472
rect 886 1468 890 1472
rect 1014 1468 1018 1472
rect 1134 1468 1138 1472
rect 1366 1468 1370 1472
rect 1382 1468 1386 1472
rect 38 1458 42 1462
rect 62 1458 66 1462
rect 110 1458 114 1462
rect 134 1458 138 1462
rect 206 1458 210 1462
rect 246 1459 250 1463
rect 366 1458 370 1462
rect 462 1458 466 1462
rect 582 1458 586 1462
rect 598 1458 602 1462
rect 646 1458 650 1462
rect 718 1458 722 1462
rect 814 1458 818 1462
rect 870 1458 874 1462
rect 950 1458 954 1462
rect 958 1458 962 1462
rect 1046 1458 1050 1462
rect 1054 1458 1058 1462
rect 1070 1458 1074 1462
rect 1094 1458 1098 1462
rect 1150 1458 1154 1462
rect 1182 1458 1186 1462
rect 1214 1458 1218 1462
rect 1246 1458 1250 1462
rect 1270 1458 1274 1462
rect 1278 1458 1282 1462
rect 1318 1458 1322 1462
rect 1350 1458 1354 1462
rect 1374 1458 1378 1462
rect 1438 1468 1442 1472
rect 1462 1468 1466 1472
rect 1494 1468 1498 1472
rect 1542 1468 1546 1472
rect 1558 1468 1562 1472
rect 1598 1468 1602 1472
rect 1646 1468 1650 1472
rect 1686 1468 1690 1472
rect 1710 1468 1714 1472
rect 1718 1468 1722 1472
rect 1734 1468 1738 1472
rect 1774 1468 1778 1472
rect 1822 1468 1826 1472
rect 1830 1468 1834 1472
rect 1846 1468 1850 1472
rect 1886 1468 1890 1472
rect 2014 1466 2018 1470
rect 2022 1468 2026 1472
rect 1486 1458 1490 1462
rect 1590 1458 1594 1462
rect 1710 1458 1714 1462
rect 1766 1458 1770 1462
rect 1798 1458 1802 1462
rect 1822 1458 1826 1462
rect 1854 1458 1858 1462
rect 1862 1458 1866 1462
rect 1886 1458 1890 1462
rect 1926 1458 1930 1462
rect 1942 1458 1946 1462
rect 1974 1458 1978 1462
rect 2046 1458 2050 1462
rect 126 1448 130 1452
rect 182 1448 186 1452
rect 190 1448 194 1452
rect 558 1448 562 1452
rect 806 1450 810 1454
rect 894 1448 898 1452
rect 1030 1448 1034 1452
rect 1062 1448 1066 1452
rect 1118 1448 1122 1452
rect 1142 1448 1146 1452
rect 1206 1448 1210 1452
rect 1238 1448 1242 1452
rect 1454 1448 1458 1452
rect 1462 1448 1466 1452
rect 1574 1448 1578 1452
rect 1638 1448 1642 1452
rect 1670 1448 1674 1452
rect 1734 1448 1738 1452
rect 1790 1448 1794 1452
rect 1934 1448 1938 1452
rect 1990 1448 1994 1452
rect 1038 1438 1042 1442
rect 1070 1438 1074 1442
rect 1078 1438 1082 1442
rect 1158 1438 1162 1442
rect 1174 1438 1178 1442
rect 1190 1438 1194 1442
rect 1222 1438 1226 1442
rect 1254 1438 1258 1442
rect 1286 1438 1290 1442
rect 1806 1438 1810 1442
rect 1862 1438 1866 1442
rect 1950 1438 1954 1442
rect 1974 1438 1978 1442
rect 310 1418 314 1422
rect 518 1418 522 1422
rect 526 1418 530 1422
rect 638 1418 642 1422
rect 678 1418 682 1422
rect 806 1418 810 1422
rect 854 1418 858 1422
rect 918 1418 922 1422
rect 1094 1418 1098 1422
rect 1166 1418 1170 1422
rect 1182 1418 1186 1422
rect 1230 1418 1234 1422
rect 1262 1418 1266 1422
rect 1278 1418 1282 1422
rect 1310 1418 1314 1422
rect 1446 1418 1450 1422
rect 1726 1418 1730 1422
rect 1782 1418 1786 1422
rect 1958 1418 1962 1422
rect 1998 1418 2002 1422
rect 2030 1418 2034 1422
rect 498 1403 502 1407
rect 505 1403 509 1407
rect 1530 1403 1534 1407
rect 1537 1403 1541 1407
rect 14 1388 18 1392
rect 158 1388 162 1392
rect 190 1388 194 1392
rect 214 1388 218 1392
rect 358 1388 362 1392
rect 1414 1388 1418 1392
rect 1454 1388 1458 1392
rect 1614 1388 1618 1392
rect 1758 1388 1762 1392
rect 1910 1388 1914 1392
rect 1926 1388 1930 1392
rect 2014 1388 2018 1392
rect 622 1368 626 1372
rect 1766 1368 1770 1372
rect 1934 1368 1938 1372
rect 158 1358 162 1362
rect 182 1358 186 1362
rect 358 1358 362 1362
rect 406 1358 410 1362
rect 446 1358 450 1362
rect 638 1358 642 1362
rect 158 1348 162 1352
rect 254 1348 258 1352
rect 342 1348 346 1352
rect 390 1348 394 1352
rect 414 1348 418 1352
rect 462 1348 466 1352
rect 502 1348 506 1352
rect 558 1348 562 1352
rect 702 1358 706 1362
rect 710 1358 714 1362
rect 782 1358 786 1362
rect 654 1348 658 1352
rect 662 1348 666 1352
rect 670 1348 674 1352
rect 734 1348 738 1352
rect 934 1358 938 1362
rect 798 1348 802 1352
rect 806 1348 810 1352
rect 886 1347 890 1351
rect 958 1348 962 1352
rect 1022 1348 1026 1352
rect 1054 1348 1058 1352
rect 1062 1348 1066 1352
rect 1086 1348 1090 1352
rect 1110 1348 1114 1352
rect 1134 1358 1138 1362
rect 1254 1358 1258 1362
rect 1294 1358 1298 1362
rect 1486 1358 1490 1362
rect 1702 1358 1706 1362
rect 1726 1358 1730 1362
rect 1782 1358 1786 1362
rect 1846 1358 1850 1362
rect 1878 1358 1882 1362
rect 1902 1358 1906 1362
rect 1950 1358 1954 1362
rect 1190 1348 1194 1352
rect 1222 1347 1226 1351
rect 1302 1348 1306 1352
rect 1318 1348 1322 1352
rect 1342 1348 1346 1352
rect 1366 1348 1370 1352
rect 1374 1348 1378 1352
rect 1398 1348 1402 1352
rect 1430 1348 1434 1352
rect 1438 1348 1442 1352
rect 1566 1348 1570 1352
rect 1614 1348 1618 1352
rect 1638 1348 1642 1352
rect 1654 1348 1658 1352
rect 1662 1348 1666 1352
rect 1686 1348 1690 1352
rect 1718 1348 1722 1352
rect 1742 1348 1746 1352
rect 1774 1348 1778 1352
rect 1790 1348 1794 1352
rect 1806 1348 1810 1352
rect 1830 1348 1834 1352
rect 1854 1348 1858 1352
rect 1862 1348 1866 1352
rect 1942 1348 1946 1352
rect 1982 1348 1986 1352
rect 110 1338 114 1342
rect 198 1338 202 1342
rect 310 1338 314 1342
rect 382 1338 386 1342
rect 422 1338 426 1342
rect 454 1338 458 1342
rect 470 1338 474 1342
rect 518 1338 522 1342
rect 622 1338 626 1342
rect 670 1338 674 1342
rect 678 1338 682 1342
rect 726 1338 730 1342
rect 742 1338 746 1342
rect 766 1338 770 1342
rect 814 1338 818 1342
rect 870 1338 874 1342
rect 918 1338 922 1342
rect 942 1338 946 1342
rect 966 1338 970 1342
rect 1046 1338 1050 1342
rect 1102 1338 1106 1342
rect 1150 1338 1154 1342
rect 1238 1338 1242 1342
rect 1270 1338 1274 1342
rect 1342 1338 1346 1342
rect 1390 1338 1394 1342
rect 1462 1338 1466 1342
rect 1526 1338 1530 1342
rect 1718 1338 1722 1342
rect 1750 1338 1754 1342
rect 1790 1338 1794 1342
rect 1806 1338 1810 1342
rect 1838 1338 1842 1342
rect 1894 1338 1898 1342
rect 1918 1338 1922 1342
rect 1958 1338 1962 1342
rect 1974 1338 1978 1342
rect 1990 1338 1994 1342
rect 2046 1338 2050 1342
rect 94 1328 98 1332
rect 294 1328 298 1332
rect 438 1328 442 1332
rect 478 1328 482 1332
rect 550 1328 554 1332
rect 758 1328 762 1332
rect 982 1328 986 1332
rect 1262 1328 1266 1332
rect 1326 1328 1330 1332
rect 1350 1328 1354 1332
rect 1614 1328 1618 1332
rect 1630 1328 1634 1332
rect 1638 1328 1642 1332
rect 1958 1328 1962 1332
rect 406 1318 410 1322
rect 430 1318 434 1322
rect 486 1318 490 1322
rect 614 1318 618 1322
rect 702 1318 706 1322
rect 718 1318 722 1322
rect 750 1318 754 1322
rect 822 1318 826 1322
rect 1070 1318 1074 1322
rect 1126 1318 1130 1322
rect 1158 1318 1162 1322
rect 1678 1318 1682 1322
rect 1702 1318 1706 1322
rect 1018 1303 1022 1307
rect 1025 1303 1029 1307
rect 254 1288 258 1292
rect 422 1288 426 1292
rect 462 1288 466 1292
rect 494 1288 498 1292
rect 726 1288 730 1292
rect 894 1288 898 1292
rect 1182 1288 1186 1292
rect 1366 1288 1370 1292
rect 1446 1288 1450 1292
rect 1694 1288 1698 1292
rect 1774 1288 1778 1292
rect 1990 1288 1994 1292
rect 2030 1288 2034 1292
rect 30 1278 34 1282
rect 110 1278 114 1282
rect 550 1278 554 1282
rect 590 1278 594 1282
rect 614 1278 618 1282
rect 870 1278 874 1282
rect 878 1278 882 1282
rect 1102 1278 1106 1282
rect 1150 1278 1154 1282
rect 1158 1278 1162 1282
rect 126 1268 130 1272
rect 174 1268 178 1272
rect 262 1268 266 1272
rect 414 1268 418 1272
rect 438 1268 442 1272
rect 470 1268 474 1272
rect 502 1268 506 1272
rect 534 1268 538 1272
rect 582 1268 586 1272
rect 606 1268 610 1272
rect 654 1268 658 1272
rect 662 1268 666 1272
rect 678 1268 682 1272
rect 694 1268 698 1272
rect 782 1268 786 1272
rect 846 1268 850 1272
rect 990 1268 994 1272
rect 1006 1268 1010 1272
rect 1054 1268 1058 1272
rect 1070 1268 1074 1272
rect 1086 1268 1090 1272
rect 1094 1268 1098 1272
rect 1238 1268 1242 1272
rect 1374 1268 1378 1272
rect 1390 1268 1394 1272
rect 1422 1268 1426 1272
rect 1542 1278 1546 1282
rect 1614 1278 1618 1282
rect 1646 1278 1650 1282
rect 1838 1278 1842 1282
rect 1998 1278 2002 1282
rect 2014 1278 2018 1282
rect 2022 1278 2026 1282
rect 1582 1268 1586 1272
rect 1598 1268 1602 1272
rect 1614 1268 1618 1272
rect 1630 1268 1634 1272
rect 54 1258 58 1262
rect 126 1258 130 1262
rect 150 1258 154 1262
rect 158 1258 162 1262
rect 198 1258 202 1262
rect 270 1258 274 1262
rect 310 1258 314 1262
rect 358 1258 362 1262
rect 374 1258 378 1262
rect 446 1258 450 1262
rect 478 1258 482 1262
rect 494 1258 498 1262
rect 518 1258 522 1262
rect 574 1258 578 1262
rect 638 1258 642 1262
rect 646 1258 650 1262
rect 670 1258 674 1262
rect 702 1258 706 1262
rect 710 1258 714 1262
rect 774 1258 778 1262
rect 838 1258 842 1262
rect 854 1258 858 1262
rect 926 1258 930 1262
rect 950 1258 954 1262
rect 1046 1258 1050 1262
rect 1078 1258 1082 1262
rect 1102 1258 1106 1262
rect 1118 1258 1122 1262
rect 1134 1258 1138 1262
rect 1174 1258 1178 1262
rect 1238 1258 1242 1262
rect 1310 1258 1314 1262
rect 1382 1258 1386 1262
rect 1478 1258 1482 1262
rect 1510 1259 1514 1263
rect 1686 1268 1690 1272
rect 1734 1268 1738 1272
rect 1790 1268 1794 1272
rect 1814 1268 1818 1272
rect 1854 1268 1858 1272
rect 1870 1268 1874 1272
rect 1894 1268 1898 1272
rect 1902 1268 1906 1272
rect 1974 1268 1978 1272
rect 1982 1268 1986 1272
rect 1574 1258 1578 1262
rect 1606 1258 1610 1262
rect 1638 1258 1642 1262
rect 1662 1258 1666 1262
rect 1670 1258 1674 1262
rect 1726 1258 1730 1262
rect 1742 1258 1746 1262
rect 1822 1258 1826 1262
rect 1918 1258 1922 1262
rect 1934 1258 1938 1262
rect 1958 1258 1962 1262
rect 2006 1258 2010 1262
rect 2046 1258 2050 1262
rect 270 1248 274 1252
rect 294 1248 298 1252
rect 430 1248 434 1252
rect 462 1248 466 1252
rect 558 1248 562 1252
rect 574 1248 578 1252
rect 590 1248 594 1252
rect 630 1248 634 1252
rect 686 1248 690 1252
rect 718 1248 722 1252
rect 822 1248 826 1252
rect 1006 1248 1010 1252
rect 1062 1248 1066 1252
rect 1406 1248 1410 1252
rect 1646 1248 1650 1252
rect 1710 1248 1714 1252
rect 1774 1248 1778 1252
rect 1798 1248 1802 1252
rect 414 1238 418 1242
rect 1198 1238 1202 1242
rect 1350 1238 1354 1242
rect 550 1228 554 1232
rect 1166 1228 1170 1232
rect 622 1218 626 1222
rect 726 1218 730 1222
rect 838 1218 842 1222
rect 862 1218 866 1222
rect 1438 1218 1442 1222
rect 1446 1218 1450 1222
rect 1758 1218 1762 1222
rect 1806 1218 1810 1222
rect 1886 1218 1890 1222
rect 1910 1218 1914 1222
rect 498 1203 502 1207
rect 505 1203 509 1207
rect 1530 1203 1534 1207
rect 1537 1203 1541 1207
rect 750 1188 754 1192
rect 790 1188 794 1192
rect 1142 1188 1146 1192
rect 1230 1188 1234 1192
rect 1630 1188 1634 1192
rect 1654 1188 1658 1192
rect 2038 1188 2042 1192
rect 646 1178 650 1182
rect 1294 1178 1298 1182
rect 1470 1179 1474 1183
rect 1710 1179 1714 1183
rect 1838 1178 1842 1182
rect 174 1168 178 1172
rect 358 1168 362 1172
rect 1622 1168 1626 1172
rect 374 1158 378 1162
rect 54 1148 58 1152
rect 142 1148 146 1152
rect 198 1148 202 1152
rect 214 1148 218 1152
rect 222 1148 226 1152
rect 246 1148 250 1152
rect 294 1148 298 1152
rect 438 1158 442 1162
rect 398 1148 402 1152
rect 422 1148 426 1152
rect 470 1148 474 1152
rect 510 1148 514 1152
rect 526 1148 530 1152
rect 534 1148 538 1152
rect 558 1158 562 1162
rect 638 1158 642 1162
rect 918 1158 922 1162
rect 1054 1158 1058 1162
rect 614 1148 618 1152
rect 622 1148 626 1152
rect 678 1148 682 1152
rect 702 1148 706 1152
rect 774 1148 778 1152
rect 870 1148 874 1152
rect 878 1148 882 1152
rect 966 1148 970 1152
rect 1190 1158 1194 1162
rect 1214 1158 1218 1162
rect 1326 1158 1330 1162
rect 1470 1156 1474 1160
rect 1518 1158 1522 1162
rect 1638 1158 1642 1162
rect 1670 1158 1674 1162
rect 1710 1156 1714 1160
rect 1078 1148 1082 1152
rect 1094 1148 1098 1152
rect 1206 1148 1210 1152
rect 1238 1148 1242 1152
rect 1246 1148 1250 1152
rect 1294 1148 1298 1152
rect 1382 1148 1386 1152
rect 1494 1148 1498 1152
rect 1510 1148 1514 1152
rect 1574 1148 1578 1152
rect 1606 1148 1610 1152
rect 1630 1148 1634 1152
rect 1654 1148 1658 1152
rect 1694 1148 1698 1152
rect 1886 1148 1890 1152
rect 1910 1148 1914 1152
rect 1974 1147 1978 1151
rect 30 1138 34 1142
rect 110 1138 114 1142
rect 270 1138 274 1142
rect 358 1138 362 1142
rect 382 1138 386 1142
rect 406 1138 410 1142
rect 414 1138 418 1142
rect 462 1138 466 1142
rect 478 1138 482 1142
rect 526 1138 530 1142
rect 582 1138 586 1142
rect 598 1138 602 1142
rect 614 1138 618 1142
rect 630 1138 634 1142
rect 742 1138 746 1142
rect 798 1138 802 1142
rect 830 1138 834 1142
rect 854 1138 858 1142
rect 862 1138 866 1142
rect 886 1138 890 1142
rect 902 1138 906 1142
rect 934 1138 938 1142
rect 1022 1138 1026 1142
rect 1062 1138 1066 1142
rect 1086 1138 1090 1142
rect 1118 1138 1122 1142
rect 1126 1138 1130 1142
rect 1174 1138 1178 1142
rect 1238 1138 1242 1142
rect 1254 1138 1258 1142
rect 1302 1138 1306 1142
rect 1310 1138 1314 1142
rect 1326 1138 1330 1142
rect 1438 1138 1442 1142
rect 1566 1138 1570 1142
rect 1598 1138 1602 1142
rect 1646 1138 1650 1142
rect 1742 1138 1746 1142
rect 238 1128 242 1132
rect 582 1128 586 1132
rect 838 1128 842 1132
rect 1270 1128 1274 1132
rect 1422 1128 1426 1132
rect 1526 1128 1530 1132
rect 1542 1128 1546 1132
rect 1582 1128 1586 1132
rect 1590 1128 1594 1132
rect 1758 1128 1762 1132
rect 94 1118 98 1122
rect 350 1118 354 1122
rect 454 1118 458 1122
rect 550 1118 554 1122
rect 590 1118 594 1122
rect 790 1118 794 1122
rect 822 1118 826 1122
rect 1022 1118 1026 1122
rect 1342 1118 1346 1122
rect 1558 1118 1562 1122
rect 1854 1118 1858 1122
rect 1018 1103 1022 1107
rect 1025 1103 1029 1107
rect 6 1088 10 1092
rect 190 1088 194 1092
rect 278 1088 282 1092
rect 446 1088 450 1092
rect 526 1088 530 1092
rect 550 1088 554 1092
rect 582 1088 586 1092
rect 670 1088 674 1092
rect 718 1088 722 1092
rect 846 1088 850 1092
rect 1270 1088 1274 1092
rect 1310 1088 1314 1092
rect 1622 1088 1626 1092
rect 1726 1088 1730 1092
rect 1990 1088 1994 1092
rect 102 1078 106 1082
rect 222 1078 226 1082
rect 270 1078 274 1082
rect 310 1078 314 1082
rect 350 1078 354 1082
rect 398 1078 402 1082
rect 454 1078 458 1082
rect 646 1078 650 1082
rect 662 1078 666 1082
rect 734 1078 738 1082
rect 782 1078 786 1082
rect 894 1078 898 1082
rect 942 1078 946 1082
rect 974 1078 978 1082
rect 1206 1078 1210 1082
rect 1382 1078 1386 1082
rect 1598 1078 1602 1082
rect 1654 1078 1658 1082
rect 1678 1078 1682 1082
rect 1686 1078 1690 1082
rect 1710 1078 1714 1082
rect 1758 1078 1762 1082
rect 62 1068 66 1072
rect 118 1068 122 1072
rect 174 1068 178 1072
rect 238 1068 242 1072
rect 294 1068 298 1072
rect 342 1068 346 1072
rect 366 1068 370 1072
rect 414 1068 418 1072
rect 438 1068 442 1072
rect 462 1068 466 1072
rect 574 1068 578 1072
rect 606 1068 610 1072
rect 614 1068 618 1072
rect 678 1068 682 1072
rect 694 1068 698 1072
rect 726 1068 730 1072
rect 854 1068 858 1072
rect 870 1068 874 1072
rect 926 1068 930 1072
rect 982 1068 986 1072
rect 1046 1068 1050 1072
rect 1134 1068 1138 1072
rect 1318 1068 1322 1072
rect 1374 1068 1378 1072
rect 1478 1068 1482 1072
rect 1614 1068 1618 1072
rect 1750 1068 1754 1072
rect 1854 1068 1858 1072
rect 1966 1068 1970 1072
rect 2014 1068 2018 1072
rect 2046 1068 2050 1072
rect 70 1059 74 1063
rect 126 1058 130 1062
rect 166 1058 170 1062
rect 174 1058 178 1062
rect 206 1058 210 1062
rect 214 1058 218 1062
rect 262 1058 266 1062
rect 286 1058 290 1062
rect 318 1058 322 1062
rect 334 1058 338 1062
rect 366 1058 370 1062
rect 382 1058 386 1062
rect 422 1058 426 1062
rect 430 1058 434 1062
rect 510 1058 514 1062
rect 566 1058 570 1062
rect 582 1058 586 1062
rect 598 1058 602 1062
rect 638 1058 642 1062
rect 686 1058 690 1062
rect 702 1058 706 1062
rect 718 1058 722 1062
rect 750 1058 754 1062
rect 798 1058 802 1062
rect 878 1058 882 1062
rect 894 1058 898 1062
rect 918 1058 922 1062
rect 958 1058 962 1062
rect 1030 1058 1034 1062
rect 1038 1058 1042 1062
rect 1110 1058 1114 1062
rect 1150 1058 1154 1062
rect 1214 1058 1218 1062
rect 1294 1058 1298 1062
rect 1326 1058 1330 1062
rect 1334 1058 1338 1062
rect 1342 1058 1346 1062
rect 1366 1058 1370 1062
rect 1454 1058 1458 1062
rect 1558 1058 1562 1062
rect 1606 1058 1610 1062
rect 1638 1058 1642 1062
rect 1662 1058 1666 1062
rect 1694 1058 1698 1062
rect 1838 1059 1842 1063
rect 1870 1058 1874 1062
rect 1878 1058 1882 1062
rect 1902 1058 1906 1062
rect 1918 1058 1922 1062
rect 1926 1058 1930 1062
rect 1958 1058 1962 1062
rect 1966 1058 1970 1062
rect 126 1048 130 1052
rect 150 1048 154 1052
rect 262 1048 266 1052
rect 854 1048 858 1052
rect 902 1048 906 1052
rect 998 1048 1002 1052
rect 1726 1048 1730 1052
rect 1942 1048 1946 1052
rect 1998 1048 2002 1052
rect 2022 1048 2026 1052
rect 1054 1038 1058 1042
rect 110 1028 114 1032
rect 1166 1028 1170 1032
rect 358 1018 362 1022
rect 654 1018 658 1022
rect 742 1018 746 1022
rect 886 1018 890 1022
rect 942 1018 946 1022
rect 966 1018 970 1022
rect 1894 1018 1898 1022
rect 2030 1018 2034 1022
rect 498 1003 502 1007
rect 505 1003 509 1007
rect 1530 1003 1534 1007
rect 1537 1003 1541 1007
rect 62 988 66 992
rect 254 988 258 992
rect 270 988 274 992
rect 486 988 490 992
rect 622 988 626 992
rect 670 988 674 992
rect 694 988 698 992
rect 902 988 906 992
rect 974 988 978 992
rect 1278 988 1282 992
rect 1822 988 1826 992
rect 302 978 306 982
rect 814 978 818 982
rect 1238 978 1242 982
rect 1134 968 1138 972
rect 1718 968 1722 972
rect 1854 968 1858 972
rect 222 958 226 962
rect 366 958 370 962
rect 398 958 402 962
rect 438 958 442 962
rect 558 958 562 962
rect 574 958 578 962
rect 766 958 770 962
rect 798 958 802 962
rect 830 958 834 962
rect 934 958 938 962
rect 1166 958 1170 962
rect 1190 958 1194 962
rect 118 948 122 952
rect 182 948 186 952
rect 190 948 194 952
rect 222 948 226 952
rect 278 948 282 952
rect 310 948 314 952
rect 342 948 346 952
rect 350 948 354 952
rect 374 948 378 952
rect 414 948 418 952
rect 430 948 434 952
rect 454 948 458 952
rect 478 948 482 952
rect 494 948 498 952
rect 558 948 562 952
rect 574 948 578 952
rect 582 948 586 952
rect 646 948 650 952
rect 654 948 658 952
rect 734 948 738 952
rect 742 948 746 952
rect 750 948 754 952
rect 758 948 762 952
rect 782 948 786 952
rect 830 948 834 952
rect 846 948 850 952
rect 870 948 874 952
rect 886 948 890 952
rect 926 948 930 952
rect 958 948 962 952
rect 990 948 994 952
rect 1022 948 1026 952
rect 1078 948 1082 952
rect 1102 948 1106 952
rect 1150 948 1154 952
rect 1470 958 1474 962
rect 1638 958 1642 962
rect 1222 948 1226 952
rect 1254 948 1258 952
rect 1262 948 1266 952
rect 1326 948 1330 952
rect 1390 948 1394 952
rect 1422 948 1426 952
rect 1454 948 1458 952
rect 1478 948 1482 952
rect 1510 948 1514 952
rect 1614 948 1618 952
rect 1678 958 1682 962
rect 1798 958 1802 962
rect 1662 948 1666 952
rect 1694 948 1698 952
rect 1718 948 1722 952
rect 1766 948 1770 952
rect 1774 948 1778 952
rect 1782 948 1786 952
rect 1806 948 1810 952
rect 1894 948 1898 952
rect 1982 948 1986 952
rect 2006 948 2010 952
rect 6 938 10 942
rect 86 938 90 942
rect 166 938 170 942
rect 174 938 178 942
rect 206 938 210 942
rect 238 938 242 942
rect 278 938 282 942
rect 318 938 322 942
rect 342 938 346 942
rect 358 938 362 942
rect 374 938 378 942
rect 422 938 426 942
rect 446 938 450 942
rect 462 938 466 942
rect 470 938 474 942
rect 510 938 514 942
rect 582 938 586 942
rect 598 938 602 942
rect 638 938 642 942
rect 718 938 722 942
rect 726 938 730 942
rect 758 938 762 942
rect 790 938 794 942
rect 822 938 826 942
rect 854 938 858 942
rect 862 938 866 942
rect 902 938 906 942
rect 918 938 922 942
rect 966 938 970 942
rect 998 938 1002 942
rect 1142 938 1146 942
rect 1158 938 1162 942
rect 1174 938 1178 942
rect 1190 938 1194 942
rect 1222 938 1226 942
rect 1302 938 1306 942
rect 1398 938 1402 942
rect 1438 938 1442 942
rect 1446 938 1450 942
rect 1486 938 1490 942
rect 1502 938 1506 942
rect 1574 938 1578 942
rect 1606 938 1610 942
rect 1614 938 1618 942
rect 1670 938 1674 942
rect 1702 938 1706 942
rect 1710 938 1714 942
rect 1758 938 1762 942
rect 1894 938 1898 942
rect 254 928 258 932
rect 262 928 266 932
rect 302 928 306 932
rect 334 928 338 932
rect 534 928 538 932
rect 614 928 618 932
rect 830 928 834 932
rect 902 928 906 932
rect 1406 928 1410 932
rect 1502 928 1506 932
rect 1526 928 1530 932
rect 1542 928 1546 932
rect 1590 928 1594 932
rect 1742 928 1746 932
rect 2014 928 2018 932
rect 62 918 66 922
rect 694 918 698 922
rect 886 918 890 922
rect 934 918 938 922
rect 974 918 978 922
rect 1382 918 1386 922
rect 1470 918 1474 922
rect 1646 918 1650 922
rect 1678 918 1682 922
rect 1934 918 1938 922
rect 1018 903 1022 907
rect 1025 903 1029 907
rect 6 888 10 892
rect 214 888 218 892
rect 494 888 498 892
rect 662 888 666 892
rect 678 888 682 892
rect 750 888 754 892
rect 838 888 842 892
rect 894 888 898 892
rect 1374 888 1378 892
rect 1574 888 1578 892
rect 1798 888 1802 892
rect 206 878 210 882
rect 374 878 378 882
rect 422 878 426 882
rect 558 878 562 882
rect 742 878 746 882
rect 934 878 938 882
rect 982 878 986 882
rect 1158 878 1162 882
rect 1286 878 1290 882
rect 1566 878 1570 882
rect 62 868 66 872
rect 86 868 90 872
rect 102 868 106 872
rect 118 868 122 872
rect 158 868 162 872
rect 174 868 178 872
rect 190 868 194 872
rect 238 868 242 872
rect 254 868 258 872
rect 294 868 298 872
rect 342 868 346 872
rect 382 868 386 872
rect 406 868 410 872
rect 438 868 442 872
rect 454 868 458 872
rect 590 868 594 872
rect 606 868 610 872
rect 638 868 642 872
rect 702 868 706 872
rect 734 868 738 872
rect 758 868 762 872
rect 806 868 810 872
rect 822 868 826 872
rect 862 868 866 872
rect 870 868 874 872
rect 918 868 922 872
rect 966 868 970 872
rect 990 868 994 872
rect 1030 868 1034 872
rect 1054 868 1058 872
rect 1062 868 1066 872
rect 1102 868 1106 872
rect 1142 868 1146 872
rect 1174 868 1178 872
rect 1270 868 1274 872
rect 1310 868 1314 872
rect 1334 868 1338 872
rect 1454 868 1458 872
rect 1494 868 1498 872
rect 1566 868 1570 872
rect 1582 868 1586 872
rect 1590 868 1594 872
rect 1710 868 1714 872
rect 1758 868 1762 872
rect 1790 868 1794 872
rect 1894 868 1898 872
rect 2014 868 2018 872
rect 2022 868 2026 872
rect 70 859 74 863
rect 142 858 146 862
rect 182 858 186 862
rect 230 858 234 862
rect 278 858 282 862
rect 358 858 362 862
rect 390 858 394 862
rect 398 858 402 862
rect 558 859 562 863
rect 630 858 634 862
rect 646 858 650 862
rect 670 858 674 862
rect 694 858 698 862
rect 734 858 738 862
rect 766 858 770 862
rect 798 858 802 862
rect 806 858 810 862
rect 854 858 858 862
rect 870 858 874 862
rect 910 858 914 862
rect 1046 858 1050 862
rect 1102 858 1106 862
rect 1166 858 1170 862
rect 1182 858 1186 862
rect 1222 858 1226 862
rect 1254 859 1258 863
rect 1302 858 1306 862
rect 1334 858 1338 862
rect 1342 858 1346 862
rect 1438 859 1442 863
rect 1486 858 1490 862
rect 1502 858 1506 862
rect 1510 858 1514 862
rect 1534 858 1538 862
rect 1590 858 1594 862
rect 1646 858 1650 862
rect 1670 858 1674 862
rect 1718 858 1722 862
rect 1766 858 1770 862
rect 1782 858 1786 862
rect 1830 858 1834 862
rect 1854 858 1858 862
rect 1902 858 1906 862
rect 1910 858 1914 862
rect 1926 858 1930 862
rect 1934 858 1938 862
rect 1942 858 1946 862
rect 2014 858 2018 862
rect 118 848 122 852
rect 158 848 162 852
rect 606 848 610 852
rect 710 848 714 852
rect 782 848 786 852
rect 830 848 834 852
rect 838 848 842 852
rect 942 848 946 852
rect 1006 848 1010 852
rect 1470 848 1474 852
rect 1718 848 1722 852
rect 1734 848 1738 852
rect 1742 848 1746 852
rect 678 838 682 842
rect 1190 838 1194 842
rect 726 828 730 832
rect 166 818 170 822
rect 662 818 666 822
rect 934 818 938 822
rect 958 818 962 822
rect 1358 818 1362 822
rect 1486 818 1490 822
rect 498 803 502 807
rect 505 803 509 807
rect 1530 803 1534 807
rect 1537 803 1541 807
rect 94 788 98 792
rect 278 788 282 792
rect 310 788 314 792
rect 726 788 730 792
rect 774 788 778 792
rect 814 788 818 792
rect 918 788 922 792
rect 1142 788 1146 792
rect 1710 788 1714 792
rect 1910 788 1914 792
rect 534 778 538 782
rect 422 768 426 772
rect 1190 768 1194 772
rect 1510 768 1514 772
rect 1814 768 1818 772
rect 1830 768 1834 772
rect 158 758 162 762
rect 302 758 306 762
rect 438 758 442 762
rect 46 748 50 752
rect 118 748 122 752
rect 126 748 130 752
rect 150 748 154 752
rect 158 748 162 752
rect 182 748 186 752
rect 214 747 218 751
rect 358 748 362 752
rect 502 758 506 762
rect 550 758 554 762
rect 678 758 682 762
rect 710 758 714 762
rect 862 758 866 762
rect 1094 758 1098 762
rect 462 748 466 752
rect 486 748 490 752
rect 494 748 498 752
rect 526 748 530 752
rect 582 748 586 752
rect 590 748 594 752
rect 622 748 626 752
rect 654 748 658 752
rect 662 748 666 752
rect 678 748 682 752
rect 694 748 698 752
rect 710 748 714 752
rect 726 748 730 752
rect 742 748 746 752
rect 766 748 770 752
rect 782 748 786 752
rect 806 748 810 752
rect 822 748 826 752
rect 838 748 842 752
rect 894 748 898 752
rect 910 748 914 752
rect 926 748 930 752
rect 958 748 962 752
rect 1022 748 1026 752
rect 1158 758 1162 762
rect 1118 748 1122 752
rect 1150 748 1154 752
rect 1158 748 1162 752
rect 1222 748 1226 752
rect 142 738 146 742
rect 182 738 186 742
rect 30 728 34 732
rect 286 738 290 742
rect 334 738 338 742
rect 366 738 370 742
rect 422 738 426 742
rect 438 738 442 742
rect 470 738 474 742
rect 478 738 482 742
rect 510 738 514 742
rect 606 738 610 742
rect 614 738 618 742
rect 630 738 634 742
rect 646 738 650 742
rect 654 738 658 742
rect 686 738 690 742
rect 1254 747 1258 751
rect 1302 748 1306 752
rect 1326 748 1330 752
rect 1358 748 1362 752
rect 1374 748 1378 752
rect 1398 758 1402 762
rect 1582 758 1586 762
rect 1614 758 1618 762
rect 1446 747 1450 751
rect 1534 748 1538 752
rect 1590 748 1594 752
rect 1598 748 1602 752
rect 1654 748 1658 752
rect 1686 748 1690 752
rect 1694 748 1698 752
rect 1734 748 1738 752
rect 1758 748 1762 752
rect 1774 748 1778 752
rect 1806 748 1810 752
rect 1846 748 1850 752
rect 1862 748 1866 752
rect 1926 748 1930 752
rect 1950 748 1954 752
rect 2006 748 2010 752
rect 718 738 722 742
rect 750 738 754 742
rect 758 738 762 742
rect 790 738 794 742
rect 798 738 802 742
rect 830 738 834 742
rect 838 738 842 742
rect 886 738 890 742
rect 902 738 906 742
rect 934 738 938 742
rect 982 738 986 742
rect 998 738 1002 742
rect 1046 738 1050 742
rect 1078 738 1082 742
rect 1126 738 1130 742
rect 1182 738 1186 742
rect 1246 738 1250 742
rect 1286 738 1290 742
rect 1350 738 1354 742
rect 1366 738 1370 742
rect 1414 738 1418 742
rect 1430 738 1434 742
rect 1542 738 1546 742
rect 1574 738 1578 742
rect 1606 738 1610 742
rect 1630 738 1634 742
rect 1678 738 1682 742
rect 1742 738 1746 742
rect 1782 738 1786 742
rect 1798 738 1802 742
rect 1934 738 1938 742
rect 2022 738 2026 742
rect 214 728 218 732
rect 246 728 250 732
rect 318 728 322 732
rect 606 728 610 732
rect 678 728 682 732
rect 942 728 946 732
rect 958 728 962 732
rect 1102 728 1106 732
rect 1134 728 1138 732
rect 1310 728 1314 732
rect 1342 728 1346 732
rect 1390 728 1394 732
rect 1550 728 1554 732
rect 1558 728 1562 732
rect 1566 728 1570 732
rect 1638 728 1642 732
rect 1726 728 1730 732
rect 1758 728 1762 732
rect 1918 728 1922 732
rect 1950 728 1954 732
rect 1974 728 1978 732
rect 294 718 298 722
rect 878 718 882 722
rect 1294 718 1298 722
rect 1614 718 1618 722
rect 1670 718 1674 722
rect 1018 703 1022 707
rect 1025 703 1029 707
rect 94 688 98 692
rect 246 688 250 692
rect 462 688 466 692
rect 582 688 586 692
rect 718 688 722 692
rect 790 688 794 692
rect 846 688 850 692
rect 878 688 882 692
rect 934 688 938 692
rect 1158 688 1162 692
rect 1398 688 1402 692
rect 1494 688 1498 692
rect 1934 688 1938 692
rect 1950 688 1954 692
rect 1990 688 1994 692
rect 2014 688 2018 692
rect 30 678 34 682
rect 366 678 370 682
rect 486 678 490 682
rect 494 678 498 682
rect 550 678 554 682
rect 694 678 698 682
rect 126 668 130 672
rect 134 668 138 672
rect 150 668 154 672
rect 166 668 170 672
rect 214 668 218 672
rect 254 668 258 672
rect 270 668 274 672
rect 286 668 290 672
rect 334 668 338 672
rect 430 668 434 672
rect 438 668 442 672
rect 478 668 482 672
rect 518 668 522 672
rect 574 668 578 672
rect 598 668 602 672
rect 614 668 618 672
rect 710 668 714 672
rect 734 678 738 682
rect 990 678 994 682
rect 1182 678 1186 682
rect 1190 678 1194 682
rect 1230 678 1234 682
rect 1294 678 1298 682
rect 1350 678 1354 682
rect 1406 678 1410 682
rect 1446 678 1450 682
rect 1502 678 1506 682
rect 1534 678 1538 682
rect 1630 678 1634 682
rect 1878 678 1882 682
rect 1982 678 1986 682
rect 2006 678 2010 682
rect 838 668 842 672
rect 870 668 874 672
rect 926 668 930 672
rect 982 668 986 672
rect 1030 668 1034 672
rect 1062 668 1066 672
rect 1174 668 1178 672
rect 1190 668 1194 672
rect 1278 668 1282 672
rect 1310 668 1314 672
rect 1326 668 1330 672
rect 1374 668 1378 672
rect 1390 668 1394 672
rect 1470 668 1474 672
rect 1478 668 1482 672
rect 1510 668 1514 672
rect 1566 668 1570 672
rect 1814 668 1818 672
rect 1870 668 1874 672
rect 1918 668 1922 672
rect 1926 668 1930 672
rect 1974 668 1978 672
rect 2022 668 2026 672
rect 46 658 50 662
rect 62 658 66 662
rect 110 658 114 662
rect 134 658 138 662
rect 190 658 194 662
rect 262 658 266 662
rect 294 658 298 662
rect 318 658 322 662
rect 366 659 370 663
rect 446 658 450 662
rect 470 658 474 662
rect 510 658 514 662
rect 566 658 570 662
rect 654 658 658 662
rect 702 658 706 662
rect 750 658 754 662
rect 758 658 762 662
rect 846 658 850 662
rect 862 658 866 662
rect 918 658 922 662
rect 1014 658 1018 662
rect 1054 658 1058 662
rect 1102 658 1106 662
rect 1126 658 1130 662
rect 1166 658 1170 662
rect 1262 659 1266 663
rect 1302 658 1306 662
rect 1326 658 1330 662
rect 1366 658 1370 662
rect 1382 658 1386 662
rect 1414 658 1418 662
rect 1446 658 1450 662
rect 1462 658 1466 662
rect 1478 658 1482 662
rect 1518 658 1522 662
rect 1582 659 1586 663
rect 1654 658 1658 662
rect 1662 658 1666 662
rect 1686 658 1690 662
rect 1694 658 1698 662
rect 1750 658 1754 662
rect 1758 658 1762 662
rect 1822 658 1826 662
rect 1846 658 1850 662
rect 1854 658 1858 662
rect 1862 658 1866 662
rect 1910 658 1914 662
rect 1918 658 1922 662
rect 1966 658 1970 662
rect 1998 658 2002 662
rect 2030 658 2034 662
rect 102 648 106 652
rect 134 648 138 652
rect 278 648 282 652
rect 310 648 314 652
rect 318 648 322 652
rect 462 648 466 652
rect 542 648 546 652
rect 550 648 554 652
rect 582 648 586 652
rect 790 648 794 652
rect 814 648 818 652
rect 846 648 850 652
rect 878 648 882 652
rect 902 648 906 652
rect 934 648 938 652
rect 958 648 962 652
rect 1022 648 1026 652
rect 1038 648 1042 652
rect 1342 648 1346 652
rect 1542 648 1546 652
rect 1678 648 1682 652
rect 1894 648 1898 652
rect 1950 648 1954 652
rect 334 638 338 642
rect 414 638 418 642
rect 526 638 530 642
rect 774 638 778 642
rect 1830 618 1834 622
rect 498 603 502 607
rect 505 603 509 607
rect 1530 603 1534 607
rect 1537 603 1541 607
rect 94 588 98 592
rect 414 588 418 592
rect 622 588 626 592
rect 870 588 874 592
rect 1070 588 1074 592
rect 1470 588 1474 592
rect 1766 588 1770 592
rect 1910 588 1914 592
rect 1926 588 1930 592
rect 758 578 762 582
rect 190 568 194 572
rect 206 568 210 572
rect 350 568 354 572
rect 526 568 530 572
rect 558 568 562 572
rect 1190 568 1194 572
rect 38 548 42 552
rect 142 548 146 552
rect 198 548 202 552
rect 230 558 234 562
rect 366 558 370 562
rect 294 548 298 552
rect 430 558 434 562
rect 382 548 386 552
rect 390 548 394 552
rect 414 548 418 552
rect 470 548 474 552
rect 558 548 562 552
rect 582 558 586 562
rect 606 558 610 562
rect 774 558 778 562
rect 622 548 626 552
rect 630 548 634 552
rect 654 548 658 552
rect 702 548 706 552
rect 774 548 778 552
rect 798 558 802 562
rect 854 558 858 562
rect 846 548 850 552
rect 870 548 874 552
rect 894 548 898 552
rect 918 558 922 562
rect 1046 558 1050 562
rect 1118 558 1122 562
rect 966 547 970 551
rect 998 548 1002 552
rect 1142 548 1146 552
rect 1158 548 1162 552
rect 1238 548 1242 552
rect 1294 548 1298 552
rect 1302 548 1306 552
rect 1318 558 1322 562
rect 1590 558 1594 562
rect 1774 558 1778 562
rect 1918 558 1922 562
rect 1998 558 2002 562
rect 1366 547 1370 551
rect 1398 548 1402 552
rect 1438 548 1442 552
rect 1502 548 1506 552
rect 1534 547 1538 551
rect 1662 547 1666 551
rect 1694 548 1698 552
rect 1702 548 1706 552
rect 1734 548 1738 552
rect 1742 548 1746 552
rect 1790 548 1794 552
rect 1830 547 1834 551
rect 1934 548 1938 552
rect 1974 548 1978 552
rect 1990 548 1994 552
rect 2046 548 2050 552
rect 110 538 114 542
rect 198 538 202 542
rect 246 538 250 542
rect 398 538 402 542
rect 406 538 410 542
rect 446 538 450 542
rect 462 538 466 542
rect 534 538 538 542
rect 550 538 554 542
rect 598 538 602 542
rect 630 538 634 542
rect 646 538 650 542
rect 710 538 714 542
rect 766 538 770 542
rect 814 538 818 542
rect 838 538 842 542
rect 878 538 882 542
rect 886 538 890 542
rect 918 538 922 542
rect 934 538 938 542
rect 1078 538 1082 542
rect 1102 538 1106 542
rect 1150 538 1154 542
rect 1166 538 1170 542
rect 1246 538 1250 542
rect 1286 538 1290 542
rect 1334 538 1338 542
rect 1350 538 1354 542
rect 1414 538 1418 542
rect 1566 538 1570 542
rect 1654 538 1658 542
rect 1750 538 1754 542
rect 1798 538 1802 542
rect 1814 538 1818 542
rect 1934 538 1938 542
rect 1942 538 1946 542
rect 2014 538 2018 542
rect 2038 538 2042 542
rect 30 528 34 532
rect 278 528 282 532
rect 662 528 666 532
rect 822 528 826 532
rect 830 528 834 532
rect 1182 528 1186 532
rect 1718 528 1722 532
rect 1990 528 1994 532
rect 2022 528 2026 532
rect 94 518 98 522
rect 1030 518 1034 522
rect 1126 518 1130 522
rect 1174 518 1178 522
rect 1454 518 1458 522
rect 1958 518 1962 522
rect 2030 518 2034 522
rect 1018 503 1022 507
rect 1025 503 1029 507
rect 62 488 66 492
rect 110 488 114 492
rect 334 488 338 492
rect 566 488 570 492
rect 590 488 594 492
rect 870 488 874 492
rect 902 488 906 492
rect 942 488 946 492
rect 1046 488 1050 492
rect 1078 488 1082 492
rect 1102 488 1106 492
rect 1166 488 1170 492
rect 1342 488 1346 492
rect 1630 488 1634 492
rect 2014 488 2018 492
rect 78 478 82 482
rect 454 478 458 482
rect 878 478 882 482
rect 910 478 914 482
rect 1054 478 1058 482
rect 1086 478 1090 482
rect 1094 478 1098 482
rect 1174 478 1178 482
rect 1246 478 1250 482
rect 1438 478 1442 482
rect 1494 478 1498 482
rect 1878 478 1882 482
rect 2030 478 2034 482
rect 6 468 10 472
rect 126 468 130 472
rect 134 468 138 472
rect 158 468 162 472
rect 190 468 194 472
rect 222 468 226 472
rect 238 468 242 472
rect 254 468 258 472
rect 278 468 282 472
rect 342 468 346 472
rect 366 468 370 472
rect 390 468 394 472
rect 510 468 514 472
rect 542 468 546 472
rect 614 468 618 472
rect 710 468 714 472
rect 822 468 826 472
rect 894 468 898 472
rect 918 468 922 472
rect 958 468 962 472
rect 974 468 978 472
rect 1006 468 1010 472
rect 1038 468 1042 472
rect 1070 468 1074 472
rect 1110 468 1114 472
rect 1118 468 1122 472
rect 1150 468 1154 472
rect 1262 468 1266 472
rect 94 458 98 462
rect 126 458 130 462
rect 174 458 178 462
rect 182 458 186 462
rect 270 459 274 463
rect 350 458 354 462
rect 422 459 426 463
rect 1302 468 1306 472
rect 1398 468 1402 472
rect 1462 468 1466 472
rect 1478 468 1482 472
rect 1518 468 1522 472
rect 1558 468 1562 472
rect 1622 468 1626 472
rect 1670 468 1674 472
rect 1678 468 1682 472
rect 1726 468 1730 472
rect 1918 468 1922 472
rect 1990 468 1994 472
rect 2006 468 2010 472
rect 2022 468 2026 472
rect 446 458 450 462
rect 518 458 522 462
rect 574 458 578 462
rect 654 458 658 462
rect 750 458 754 462
rect 806 458 810 462
rect 822 458 826 462
rect 846 458 850 462
rect 854 458 858 462
rect 862 458 866 462
rect 886 458 890 462
rect 926 458 930 462
rect 966 458 970 462
rect 982 458 986 462
rect 1030 458 1034 462
rect 1062 458 1066 462
rect 1118 458 1122 462
rect 1142 458 1146 462
rect 1158 458 1162 462
rect 1222 458 1226 462
rect 1278 458 1282 462
rect 1294 458 1298 462
rect 1334 458 1338 462
rect 1406 459 1410 463
rect 1454 458 1458 462
rect 1486 458 1490 462
rect 1510 458 1514 462
rect 1558 458 1562 462
rect 1574 458 1578 462
rect 1598 458 1602 462
rect 1614 458 1618 462
rect 1670 458 1674 462
rect 1782 458 1786 462
rect 1806 458 1810 462
rect 1854 458 1858 462
rect 1862 458 1866 462
rect 1870 458 1874 462
rect 1902 458 1906 462
rect 1958 458 1962 462
rect 2046 458 2050 462
rect 150 448 154 452
rect 222 448 226 452
rect 374 448 378 452
rect 534 448 538 452
rect 566 448 570 452
rect 942 448 946 452
rect 950 448 954 452
rect 1126 448 1130 452
rect 1278 448 1282 452
rect 1494 448 1498 452
rect 1646 448 1650 452
rect 1702 448 1706 452
rect 1982 438 1986 442
rect 694 418 698 422
rect 1318 418 1322 422
rect 1550 418 1554 422
rect 1590 418 1594 422
rect 1686 418 1690 422
rect 1710 418 1714 422
rect 1734 418 1738 422
rect 498 403 502 407
rect 505 403 509 407
rect 1530 403 1534 407
rect 1537 403 1541 407
rect 110 388 114 392
rect 438 388 442 392
rect 534 388 538 392
rect 550 388 554 392
rect 582 388 586 392
rect 750 388 754 392
rect 798 388 802 392
rect 894 388 898 392
rect 1046 388 1050 392
rect 1486 388 1490 392
rect 1566 388 1570 392
rect 1950 388 1954 392
rect 318 368 322 372
rect 1086 368 1090 372
rect 1374 368 1378 372
rect 1398 368 1402 372
rect 374 358 378 362
rect 454 358 458 362
rect 590 358 594 362
rect 630 358 634 362
rect 6 348 10 352
rect 54 348 58 352
rect 126 348 130 352
rect 150 348 154 352
rect 158 348 162 352
rect 182 348 186 352
rect 190 348 194 352
rect 222 348 226 352
rect 270 348 274 352
rect 334 348 338 352
rect 342 348 346 352
rect 398 348 402 352
rect 438 348 442 352
rect 462 348 466 352
rect 478 348 482 352
rect 510 348 514 352
rect 558 348 562 352
rect 614 348 618 352
rect 646 348 650 352
rect 662 348 666 352
rect 670 348 674 352
rect 686 358 690 362
rect 806 358 810 362
rect 734 348 738 352
rect 798 348 802 352
rect 814 348 818 352
rect 822 348 826 352
rect 846 348 850 352
rect 870 358 874 362
rect 1790 358 1794 362
rect 934 348 938 352
rect 990 348 994 352
rect 1038 348 1042 352
rect 1054 348 1058 352
rect 1078 348 1082 352
rect 1102 348 1106 352
rect 1110 348 1114 352
rect 1118 348 1122 352
rect 1206 348 1210 352
rect 1278 348 1282 352
rect 1326 348 1330 352
rect 1334 348 1338 352
rect 1350 348 1354 352
rect 1358 348 1362 352
rect 1422 348 1426 352
rect 1622 348 1626 352
rect 1694 348 1698 352
rect 1726 348 1730 352
rect 1734 348 1738 352
rect 1742 348 1746 352
rect 1766 348 1770 352
rect 1814 348 1818 352
rect 1846 348 1850 352
rect 1886 348 1890 352
rect 1894 348 1898 352
rect 1982 348 1986 352
rect 2014 347 2018 351
rect 30 338 34 342
rect 62 338 66 342
rect 166 338 170 342
rect 326 338 330 342
rect 358 338 362 342
rect 406 338 410 342
rect 430 338 434 342
rect 470 338 474 342
rect 518 338 522 342
rect 614 338 618 342
rect 622 338 626 342
rect 654 338 658 342
rect 702 338 706 342
rect 774 338 778 342
rect 830 338 834 342
rect 838 338 842 342
rect 862 338 866 342
rect 974 338 978 342
rect 1062 338 1066 342
rect 1126 338 1130 342
rect 1158 338 1162 342
rect 1246 338 1250 342
rect 1302 338 1306 342
rect 1462 338 1466 342
rect 1550 338 1554 342
rect 1662 338 1666 342
rect 1718 338 1722 342
rect 1774 338 1778 342
rect 1838 338 1842 342
rect 1846 338 1850 342
rect 6 328 10 332
rect 166 328 170 332
rect 254 328 258 332
rect 382 328 386 332
rect 422 328 426 332
rect 486 328 490 332
rect 534 328 538 332
rect 542 328 546 332
rect 566 328 570 332
rect 582 328 586 332
rect 782 328 786 332
rect 1006 328 1010 332
rect 1142 328 1146 332
rect 1262 328 1266 332
rect 1678 328 1682 332
rect 1790 328 1794 332
rect 1798 328 1802 332
rect 134 318 138 322
rect 206 318 210 322
rect 390 318 394 322
rect 414 318 418 322
rect 718 318 722 322
rect 1134 318 1138 322
rect 1294 318 1298 322
rect 1710 318 1714 322
rect 1830 318 1834 322
rect 1018 303 1022 307
rect 1025 303 1029 307
rect 6 288 10 292
rect 102 288 106 292
rect 286 288 290 292
rect 438 288 442 292
rect 590 288 594 292
rect 694 288 698 292
rect 750 288 754 292
rect 862 288 866 292
rect 1054 288 1058 292
rect 1278 288 1282 292
rect 1430 288 1434 292
rect 1446 288 1450 292
rect 1574 288 1578 292
rect 1646 288 1650 292
rect 1678 288 1682 292
rect 1918 288 1922 292
rect 318 278 322 282
rect 614 278 618 282
rect 1046 278 1050 282
rect 62 268 66 272
rect 206 268 210 272
rect 254 268 258 272
rect 342 268 346 272
rect 358 268 362 272
rect 446 268 450 272
rect 494 268 498 272
rect 502 268 506 272
rect 550 268 554 272
rect 598 268 602 272
rect 630 268 634 272
rect 662 268 666 272
rect 670 268 674 272
rect 726 268 730 272
rect 782 268 786 272
rect 830 268 834 272
rect 838 268 842 272
rect 918 268 922 272
rect 934 268 938 272
rect 950 268 954 272
rect 1062 268 1066 272
rect 1422 278 1426 282
rect 1118 268 1122 272
rect 1126 268 1130 272
rect 1158 268 1162 272
rect 1190 268 1194 272
rect 1222 268 1226 272
rect 1246 268 1250 272
rect 1270 268 1274 272
rect 1318 268 1322 272
rect 1326 268 1330 272
rect 1406 268 1410 272
rect 1566 268 1570 272
rect 1590 278 1594 282
rect 1614 278 1618 282
rect 1790 278 1794 282
rect 1934 278 1938 282
rect 1942 278 1946 282
rect 1630 268 1634 272
rect 1670 268 1674 272
rect 1758 268 1762 272
rect 1926 268 1930 272
rect 70 259 74 263
rect 134 258 138 262
rect 166 259 170 263
rect 230 258 234 262
rect 334 258 338 262
rect 382 258 386 262
rect 454 258 458 262
rect 542 258 546 262
rect 558 258 562 262
rect 606 258 610 262
rect 630 258 634 262
rect 662 258 666 262
rect 678 258 682 262
rect 726 258 730 262
rect 742 258 746 262
rect 766 258 770 262
rect 774 258 778 262
rect 814 258 818 262
rect 822 258 826 262
rect 830 258 834 262
rect 870 258 874 262
rect 878 258 882 262
rect 902 258 906 262
rect 926 258 930 262
rect 958 258 962 262
rect 974 258 978 262
rect 982 258 986 262
rect 990 258 994 262
rect 1014 258 1018 262
rect 1070 258 1074 262
rect 1094 258 1098 262
rect 1126 258 1130 262
rect 1150 258 1154 262
rect 1190 258 1194 262
rect 1198 258 1202 262
rect 1214 258 1218 262
rect 1238 258 1242 262
rect 1262 258 1266 262
rect 1310 258 1314 262
rect 1366 258 1370 262
rect 1438 258 1442 262
rect 1486 258 1490 262
rect 1510 259 1514 263
rect 1542 258 1546 262
rect 1558 258 1562 262
rect 1606 258 1610 262
rect 1622 258 1626 262
rect 1638 258 1642 262
rect 1670 258 1674 262
rect 1718 258 1722 262
rect 1806 258 1810 262
rect 1830 258 1834 262
rect 1870 258 1874 262
rect 1878 258 1882 262
rect 1902 258 1906 262
rect 1942 258 1946 262
rect 1958 258 1962 262
rect 1982 258 1986 262
rect 2014 258 2018 262
rect 2022 258 2026 262
rect 310 248 314 252
rect 454 248 458 252
rect 478 248 482 252
rect 574 248 578 252
rect 638 248 642 252
rect 654 248 658 252
rect 694 248 698 252
rect 702 248 706 252
rect 718 248 722 252
rect 798 248 802 252
rect 862 248 866 252
rect 942 248 946 252
rect 974 248 978 252
rect 1134 248 1138 252
rect 1166 248 1170 252
rect 1198 248 1202 252
rect 1254 248 1258 252
rect 1294 248 1298 252
rect 1646 248 1650 252
rect 1462 238 1466 242
rect 1694 238 1698 242
rect 894 218 898 222
rect 1006 218 1010 222
rect 1102 218 1106 222
rect 1182 218 1186 222
rect 1894 218 1898 222
rect 1966 218 1970 222
rect 1998 218 2002 222
rect 2046 218 2050 222
rect 498 203 502 207
rect 505 203 509 207
rect 1530 203 1534 207
rect 1537 203 1541 207
rect 374 188 378 192
rect 590 188 594 192
rect 622 188 626 192
rect 798 188 802 192
rect 830 188 834 192
rect 990 188 994 192
rect 1046 188 1050 192
rect 1302 188 1306 192
rect 1966 188 1970 192
rect 1998 188 2002 192
rect 494 178 498 182
rect 1470 178 1474 182
rect 246 168 250 172
rect 1486 168 1490 172
rect 54 148 58 152
rect 62 148 66 152
rect 102 148 106 152
rect 134 148 138 152
rect 190 148 194 152
rect 206 148 210 152
rect 262 148 266 152
rect 270 148 274 152
rect 286 158 290 162
rect 318 148 322 152
rect 342 158 346 162
rect 398 158 402 162
rect 382 148 386 152
rect 438 148 442 152
rect 526 148 530 152
rect 534 148 538 152
rect 550 158 554 162
rect 742 158 746 162
rect 774 158 778 162
rect 854 158 858 162
rect 598 148 602 152
rect 102 138 106 142
rect 110 138 114 142
rect 254 138 258 142
rect 302 138 306 142
rect 310 138 314 142
rect 358 138 362 142
rect 686 147 690 151
rect 726 148 730 152
rect 758 148 762 152
rect 790 148 794 152
rect 814 148 818 152
rect 1158 158 1162 162
rect 878 148 882 152
rect 942 148 946 152
rect 1022 148 1026 152
rect 1102 148 1106 152
rect 1174 148 1178 152
rect 1182 148 1186 152
rect 1222 147 1226 151
rect 1366 148 1370 152
rect 1374 148 1378 152
rect 1414 148 1418 152
rect 1430 148 1434 152
rect 1462 148 1466 152
rect 1502 148 1506 152
rect 1510 148 1514 152
rect 1598 148 1602 152
rect 1630 148 1634 152
rect 1654 148 1658 152
rect 1686 148 1690 152
rect 1758 148 1762 152
rect 1782 148 1786 152
rect 1814 148 1818 152
rect 1838 148 1842 152
rect 1870 148 1874 152
rect 1902 147 1906 151
rect 1974 148 1978 152
rect 2006 148 2010 152
rect 438 138 442 142
rect 518 138 522 142
rect 566 138 570 142
rect 614 138 618 142
rect 702 138 706 142
rect 718 138 722 142
rect 750 138 754 142
rect 814 138 818 142
rect 838 138 842 142
rect 886 138 890 142
rect 998 138 1002 142
rect 1102 138 1106 142
rect 1142 138 1146 142
rect 1190 138 1194 142
rect 1206 138 1210 142
rect 1358 138 1362 142
rect 1454 138 1458 142
rect 1622 138 1626 142
rect 1678 138 1682 142
rect 1694 138 1698 142
rect 1806 138 1810 142
rect 1862 138 1866 142
rect 1886 138 1890 142
rect 118 128 122 132
rect 150 128 154 132
rect 366 128 370 132
rect 574 128 578 132
rect 614 128 618 132
rect 822 128 826 132
rect 918 128 922 132
rect 982 128 986 132
rect 998 128 1002 132
rect 1006 128 1010 132
rect 1254 128 1258 132
rect 1414 128 1418 132
rect 1446 128 1450 132
rect 1566 128 1570 132
rect 1638 128 1642 132
rect 1766 128 1770 132
rect 1822 128 1826 132
rect 2006 128 2010 132
rect 334 118 338 122
rect 398 118 402 122
rect 742 118 746 122
rect 862 118 866 122
rect 1390 118 1394 122
rect 1614 118 1618 122
rect 1670 118 1674 122
rect 1798 118 1802 122
rect 1854 118 1858 122
rect 1990 118 1994 122
rect 2038 118 2042 122
rect 1018 103 1022 107
rect 1025 103 1029 107
rect 62 88 66 92
rect 390 88 394 92
rect 430 88 434 92
rect 782 88 786 92
rect 790 88 794 92
rect 910 88 914 92
rect 1022 88 1026 92
rect 1230 88 1234 92
rect 1326 88 1330 92
rect 1526 88 1530 92
rect 1630 88 1634 92
rect 1638 88 1642 92
rect 1734 88 1738 92
rect 1830 88 1834 92
rect 2030 88 2034 92
rect 246 78 250 82
rect 598 78 602 82
rect 614 78 618 82
rect 1190 78 1194 82
rect 6 68 10 72
rect 78 68 82 72
rect 142 68 146 72
rect 158 68 162 72
rect 270 68 274 72
rect 286 68 290 72
rect 310 68 314 72
rect 422 68 426 72
rect 654 68 658 72
rect 686 68 690 72
rect 702 68 706 72
rect 806 68 810 72
rect 822 68 826 72
rect 1102 68 1106 72
rect 1118 68 1122 72
rect 1134 68 1138 72
rect 1166 68 1170 72
rect 1374 78 1378 82
rect 1406 78 1410 82
rect 1622 78 1626 82
rect 1214 68 1218 72
rect 1310 68 1314 72
rect 1438 68 1442 72
rect 1502 68 1506 72
rect 1606 68 1610 72
rect 1718 68 1722 72
rect 1886 68 1890 72
rect 2006 68 2010 72
rect 2022 68 2026 72
rect 182 58 186 62
rect 262 58 266 62
rect 294 58 298 62
rect 334 58 338 62
rect 414 58 418 62
rect 462 58 466 62
rect 486 58 490 62
rect 574 58 578 62
rect 678 58 682 62
rect 742 58 746 62
rect 846 58 850 62
rect 870 58 874 62
rect 942 58 946 62
rect 966 58 970 62
rect 1054 58 1058 62
rect 1086 59 1090 63
rect 1158 58 1162 62
rect 1174 58 1178 62
rect 1206 58 1210 62
rect 1222 58 1226 62
rect 1270 58 1274 62
rect 1390 58 1394 62
rect 1590 59 1594 63
rect 1678 58 1682 62
rect 1766 58 1770 62
rect 1798 59 1802 63
rect 1862 58 1866 62
rect 1870 58 1874 62
rect 1958 58 1962 62
rect 398 48 402 52
rect 414 48 418 52
rect 654 48 658 52
rect 790 48 794 52
rect 1134 48 1138 52
rect 498 3 502 7
rect 505 3 509 7
rect 1530 3 1534 7
rect 1537 3 1541 7
<< metal2 >>
rect 118 1828 122 1832
rect 830 1828 834 1832
rect 1934 1828 1938 1832
rect 1958 1828 1962 1832
rect 118 1792 121 1828
rect 496 1803 498 1807
rect 502 1803 505 1807
rect 509 1803 512 1807
rect 830 1802 833 1828
rect 1528 1803 1530 1807
rect 1534 1803 1537 1807
rect 1541 1803 1544 1807
rect 174 1792 177 1798
rect 10 1788 14 1791
rect 30 1782 33 1788
rect 22 1691 25 1748
rect 18 1688 25 1691
rect 6 1572 9 1578
rect 30 1552 33 1568
rect 46 1562 49 1748
rect 54 1742 57 1788
rect 350 1762 353 1788
rect 598 1762 601 1788
rect 126 1742 129 1758
rect 674 1748 678 1751
rect 54 1592 57 1738
rect 94 1682 97 1688
rect 110 1682 113 1718
rect 142 1702 145 1748
rect 150 1742 153 1748
rect 166 1692 169 1748
rect 190 1692 193 1698
rect 286 1682 289 1728
rect 302 1702 305 1738
rect 42 1548 46 1551
rect 22 1501 25 1548
rect 94 1542 97 1678
rect 14 1498 25 1501
rect 14 1392 17 1498
rect 30 1332 33 1468
rect 38 1462 41 1468
rect 62 1462 65 1538
rect 102 1492 105 1548
rect 110 1512 113 1668
rect 230 1662 233 1668
rect 162 1658 166 1661
rect 158 1622 161 1648
rect 270 1621 273 1678
rect 286 1642 289 1668
rect 334 1662 337 1748
rect 350 1742 353 1748
rect 374 1742 377 1748
rect 362 1688 366 1691
rect 398 1672 401 1748
rect 406 1722 409 1728
rect 446 1682 449 1718
rect 494 1712 497 1748
rect 534 1722 537 1728
rect 262 1618 273 1621
rect 318 1622 321 1650
rect 178 1548 181 1551
rect 166 1532 169 1548
rect 94 1482 97 1488
rect 134 1472 137 1528
rect 150 1502 153 1528
rect 146 1488 150 1491
rect 158 1482 161 1518
rect 166 1472 169 1478
rect 214 1472 217 1548
rect 262 1532 265 1618
rect 326 1562 329 1588
rect 334 1552 337 1658
rect 350 1552 353 1648
rect 438 1552 441 1558
rect 262 1482 265 1528
rect 278 1492 281 1538
rect 334 1501 337 1548
rect 334 1498 345 1501
rect 114 1468 118 1471
rect 178 1468 182 1471
rect 194 1468 198 1471
rect 102 1442 105 1468
rect 114 1458 118 1461
rect 126 1452 129 1468
rect 134 1452 137 1458
rect 94 1332 97 1338
rect 30 1282 33 1328
rect 110 1312 113 1338
rect 110 1282 113 1288
rect 30 1142 33 1278
rect 122 1268 126 1271
rect 54 1262 57 1268
rect 130 1258 134 1261
rect 54 1092 57 1148
rect 110 1142 113 1148
rect 94 1091 97 1118
rect 94 1088 105 1091
rect 6 1082 9 1088
rect 102 1082 105 1088
rect 126 1072 129 1258
rect 142 1161 145 1458
rect 182 1452 185 1458
rect 190 1392 193 1448
rect 206 1442 209 1458
rect 214 1452 217 1468
rect 158 1362 161 1388
rect 182 1352 185 1358
rect 158 1342 161 1348
rect 198 1342 201 1418
rect 210 1388 214 1391
rect 150 1282 153 1298
rect 198 1282 201 1338
rect 230 1332 233 1468
rect 246 1463 249 1468
rect 306 1418 310 1421
rect 342 1352 345 1498
rect 254 1342 257 1348
rect 294 1322 297 1328
rect 150 1262 153 1278
rect 254 1272 257 1288
rect 158 1252 161 1258
rect 174 1172 177 1268
rect 262 1262 265 1268
rect 270 1262 273 1288
rect 198 1252 201 1258
rect 142 1158 153 1161
rect 142 1132 145 1148
rect 122 1068 126 1071
rect 62 992 65 1068
rect 150 1062 153 1158
rect 214 1152 217 1258
rect 222 1152 225 1158
rect 246 1152 249 1258
rect 274 1248 278 1251
rect 202 1148 206 1151
rect 166 1062 169 1098
rect 186 1088 190 1091
rect 174 1072 177 1078
rect 214 1062 217 1148
rect 270 1142 273 1148
rect 234 1128 238 1131
rect 222 1082 225 1088
rect 278 1082 281 1088
rect 266 1078 270 1081
rect 242 1068 246 1071
rect 70 1052 73 1059
rect 130 1058 134 1061
rect 150 1052 153 1058
rect 126 1042 129 1048
rect 110 1032 113 1038
rect 6 942 9 988
rect 122 948 126 951
rect 6 882 9 888
rect 62 872 65 918
rect 86 872 89 938
rect 150 902 153 1048
rect 174 942 177 1058
rect 206 1032 209 1058
rect 214 1052 217 1058
rect 226 958 230 961
rect 182 952 185 958
rect 194 948 198 951
rect 206 942 209 948
rect 162 938 166 941
rect 174 892 177 938
rect 102 872 105 878
rect 70 863 73 868
rect 118 862 121 868
rect 94 792 97 818
rect 118 812 121 848
rect 142 812 145 858
rect 150 752 153 888
rect 158 862 161 868
rect 174 862 177 868
rect 182 862 185 878
rect 190 872 193 878
rect 158 832 161 848
rect 166 761 169 818
rect 162 758 169 761
rect 182 752 185 828
rect 50 748 54 751
rect 130 748 134 751
rect 162 748 166 751
rect 118 742 121 748
rect 142 742 145 748
rect 30 682 33 728
rect 150 712 153 748
rect 182 732 185 738
rect 98 688 102 691
rect 150 672 153 688
rect 138 668 142 671
rect 50 658 54 661
rect 62 652 65 658
rect 102 652 105 668
rect 114 658 118 661
rect 30 532 33 538
rect 10 468 14 471
rect 10 348 14 351
rect 30 342 33 528
rect 38 512 41 548
rect 62 492 65 648
rect 126 641 129 668
rect 134 652 137 658
rect 126 638 137 641
rect 94 592 97 608
rect 110 532 113 538
rect 90 518 94 521
rect 78 482 81 518
rect 110 492 113 508
rect 126 472 129 588
rect 134 542 137 638
rect 142 552 145 568
rect 94 462 97 468
rect 122 458 126 461
rect 114 388 118 391
rect 54 352 57 368
rect 126 352 129 458
rect 134 392 137 468
rect 150 462 153 658
rect 166 652 169 668
rect 182 662 185 728
rect 190 662 193 678
rect 150 452 153 458
rect 158 372 161 468
rect 182 462 185 558
rect 190 552 193 568
rect 198 562 201 898
rect 206 882 209 918
rect 214 892 217 908
rect 222 862 225 948
rect 238 942 241 1068
rect 286 1062 289 1278
rect 294 1252 297 1288
rect 310 1282 313 1338
rect 310 1262 313 1268
rect 350 1262 353 1548
rect 358 1532 361 1538
rect 382 1532 385 1548
rect 446 1542 449 1678
rect 462 1632 465 1668
rect 510 1662 513 1708
rect 534 1662 537 1668
rect 514 1658 518 1661
rect 494 1631 497 1650
rect 496 1603 498 1607
rect 502 1603 505 1607
rect 509 1603 512 1607
rect 550 1602 553 1738
rect 574 1672 577 1708
rect 606 1692 609 1748
rect 774 1742 777 1748
rect 798 1742 801 1748
rect 814 1742 817 1798
rect 918 1752 921 1788
rect 958 1760 961 1779
rect 1454 1762 1457 1788
rect 1510 1762 1513 1788
rect 1758 1762 1761 1788
rect 1934 1762 1937 1828
rect 1950 1762 1953 1768
rect 1934 1752 1937 1758
rect 918 1742 921 1748
rect 942 1742 945 1748
rect 850 1738 854 1741
rect 626 1718 633 1721
rect 630 1672 633 1718
rect 654 1692 657 1738
rect 662 1732 665 1738
rect 574 1662 577 1668
rect 582 1652 585 1668
rect 590 1622 593 1658
rect 614 1622 617 1648
rect 526 1562 529 1568
rect 522 1548 526 1551
rect 358 1472 361 1478
rect 366 1462 369 1518
rect 398 1472 401 1528
rect 446 1472 449 1538
rect 494 1482 497 1518
rect 358 1362 361 1388
rect 382 1342 385 1358
rect 390 1292 393 1348
rect 362 1258 366 1261
rect 374 1252 377 1258
rect 398 1182 401 1468
rect 462 1462 465 1468
rect 518 1462 521 1538
rect 550 1482 553 1538
rect 558 1502 561 1618
rect 630 1592 633 1668
rect 646 1662 649 1668
rect 570 1558 574 1561
rect 570 1548 574 1551
rect 538 1478 542 1481
rect 574 1472 577 1548
rect 598 1542 601 1548
rect 586 1538 590 1541
rect 598 1522 601 1528
rect 614 1492 617 1558
rect 630 1551 633 1558
rect 630 1482 633 1488
rect 638 1472 641 1658
rect 646 1542 649 1658
rect 662 1552 665 1728
rect 686 1682 689 1718
rect 674 1658 678 1661
rect 562 1468 566 1471
rect 586 1468 590 1471
rect 542 1452 545 1468
rect 518 1422 521 1448
rect 558 1432 561 1448
rect 582 1432 585 1458
rect 590 1442 593 1468
rect 646 1462 649 1538
rect 654 1492 657 1518
rect 662 1482 665 1548
rect 670 1482 673 1508
rect 598 1452 601 1458
rect 496 1403 498 1407
rect 502 1403 505 1407
rect 509 1403 512 1407
rect 406 1332 409 1358
rect 418 1348 422 1351
rect 418 1338 422 1341
rect 406 1262 409 1318
rect 422 1292 425 1328
rect 430 1312 433 1318
rect 438 1292 441 1328
rect 446 1322 449 1358
rect 462 1352 465 1368
rect 498 1348 502 1351
rect 470 1342 473 1348
rect 518 1342 521 1418
rect 526 1372 529 1418
rect 562 1348 566 1351
rect 454 1332 457 1338
rect 446 1312 449 1318
rect 414 1242 417 1268
rect 430 1252 433 1288
rect 438 1272 441 1278
rect 298 1148 302 1151
rect 358 1142 361 1168
rect 374 1132 377 1158
rect 414 1152 417 1238
rect 430 1172 433 1248
rect 438 1222 441 1268
rect 446 1262 449 1298
rect 458 1288 462 1291
rect 470 1282 473 1338
rect 478 1332 481 1338
rect 486 1272 489 1318
rect 494 1292 497 1298
rect 502 1272 505 1278
rect 474 1268 478 1271
rect 514 1258 518 1261
rect 462 1242 465 1248
rect 478 1232 481 1258
rect 494 1232 497 1258
rect 422 1152 425 1158
rect 438 1152 441 1158
rect 382 1142 385 1148
rect 350 1082 353 1118
rect 398 1102 401 1148
rect 418 1138 422 1141
rect 406 1132 409 1138
rect 446 1092 449 1228
rect 462 1142 465 1178
rect 470 1152 473 1218
rect 496 1203 498 1207
rect 502 1203 505 1207
rect 509 1203 512 1207
rect 526 1152 529 1318
rect 550 1311 553 1328
rect 542 1308 553 1311
rect 558 1312 561 1328
rect 598 1322 601 1448
rect 638 1371 641 1418
rect 638 1368 649 1371
rect 622 1342 625 1368
rect 638 1342 641 1358
rect 534 1242 537 1268
rect 542 1252 545 1308
rect 558 1281 561 1308
rect 554 1278 561 1281
rect 574 1262 577 1288
rect 614 1282 617 1318
rect 594 1278 598 1281
rect 606 1272 609 1278
rect 586 1268 590 1271
rect 646 1262 649 1368
rect 654 1352 657 1358
rect 662 1352 665 1358
rect 670 1352 673 1478
rect 678 1412 681 1418
rect 686 1362 689 1678
rect 702 1672 705 1738
rect 714 1718 718 1721
rect 750 1662 753 1738
rect 822 1712 825 1718
rect 794 1668 801 1671
rect 818 1668 822 1671
rect 710 1562 713 1618
rect 710 1552 713 1558
rect 718 1552 721 1659
rect 790 1652 793 1658
rect 798 1622 801 1668
rect 822 1622 825 1648
rect 838 1642 841 1668
rect 902 1662 905 1668
rect 910 1651 913 1738
rect 926 1672 929 1728
rect 990 1692 993 1738
rect 1006 1732 1009 1738
rect 1016 1703 1018 1707
rect 1022 1703 1025 1707
rect 1029 1703 1032 1707
rect 970 1688 974 1691
rect 1094 1682 1097 1728
rect 1118 1722 1121 1748
rect 1142 1742 1145 1748
rect 1214 1742 1217 1748
rect 1350 1742 1353 1748
rect 1462 1742 1465 1748
rect 1510 1742 1513 1748
rect 1150 1732 1153 1738
rect 1294 1732 1297 1738
rect 1390 1732 1393 1738
rect 1226 1728 1230 1731
rect 990 1672 993 1678
rect 1006 1672 1009 1678
rect 1046 1672 1049 1678
rect 1038 1668 1046 1671
rect 1178 1668 1182 1671
rect 902 1648 913 1651
rect 942 1652 945 1668
rect 738 1558 742 1561
rect 750 1542 753 1608
rect 758 1572 761 1618
rect 782 1612 785 1618
rect 838 1592 841 1638
rect 758 1542 761 1568
rect 774 1562 777 1568
rect 798 1562 801 1588
rect 770 1538 774 1541
rect 694 1512 697 1518
rect 702 1382 705 1538
rect 750 1512 753 1538
rect 718 1462 721 1498
rect 758 1482 761 1488
rect 702 1352 705 1358
rect 710 1342 713 1358
rect 734 1352 737 1358
rect 774 1352 777 1468
rect 814 1462 817 1548
rect 846 1542 849 1548
rect 862 1532 865 1638
rect 902 1552 905 1648
rect 974 1572 977 1578
rect 958 1542 961 1558
rect 982 1542 985 1638
rect 990 1552 993 1658
rect 1030 1612 1033 1618
rect 1038 1592 1041 1668
rect 1006 1532 1009 1538
rect 1046 1532 1049 1538
rect 862 1492 865 1528
rect 842 1478 846 1481
rect 890 1468 894 1471
rect 806 1422 809 1450
rect 782 1362 785 1398
rect 806 1352 809 1398
rect 794 1348 798 1351
rect 742 1342 745 1348
rect 666 1338 670 1341
rect 678 1322 681 1338
rect 678 1272 681 1278
rect 694 1272 697 1338
rect 702 1292 705 1318
rect 666 1268 670 1271
rect 578 1248 590 1251
rect 558 1242 561 1248
rect 630 1232 633 1248
rect 550 1222 553 1228
rect 534 1152 537 1158
rect 470 1142 473 1148
rect 482 1138 486 1141
rect 454 1112 457 1118
rect 470 1102 473 1138
rect 478 1132 481 1138
rect 314 1078 318 1081
rect 298 1068 302 1071
rect 346 1068 350 1071
rect 266 1058 270 1061
rect 322 1058 326 1061
rect 358 1061 361 1088
rect 470 1082 473 1098
rect 402 1078 406 1081
rect 458 1078 462 1081
rect 438 1072 441 1078
rect 510 1072 513 1148
rect 558 1142 561 1158
rect 582 1142 585 1178
rect 614 1152 617 1188
rect 622 1152 625 1218
rect 638 1192 641 1258
rect 654 1242 657 1268
rect 702 1262 705 1268
rect 666 1258 670 1261
rect 710 1252 713 1258
rect 718 1252 721 1318
rect 726 1292 729 1338
rect 642 1178 646 1181
rect 642 1158 649 1161
rect 522 1138 526 1141
rect 602 1138 606 1141
rect 634 1138 638 1141
rect 614 1132 617 1138
rect 526 1092 529 1128
rect 550 1112 553 1118
rect 582 1102 585 1128
rect 550 1092 553 1098
rect 578 1088 582 1091
rect 370 1068 374 1071
rect 418 1068 422 1071
rect 458 1068 462 1071
rect 574 1062 577 1068
rect 358 1058 366 1061
rect 514 1058 518 1061
rect 590 1061 593 1118
rect 590 1058 598 1061
rect 254 1048 262 1051
rect 254 992 257 1048
rect 334 1042 337 1058
rect 270 992 273 1038
rect 278 952 281 988
rect 302 972 305 978
rect 338 948 342 951
rect 358 951 361 1018
rect 366 962 369 968
rect 354 948 361 951
rect 374 952 377 1028
rect 382 992 385 1058
rect 422 1052 425 1058
rect 430 1052 433 1058
rect 398 962 401 1038
rect 496 1003 498 1007
rect 502 1003 505 1007
rect 509 1003 512 1007
rect 482 988 486 991
rect 230 938 238 941
rect 230 882 233 938
rect 266 928 270 931
rect 254 892 257 928
rect 278 912 281 938
rect 230 862 233 878
rect 254 872 257 878
rect 222 792 225 858
rect 238 802 241 868
rect 278 862 281 878
rect 274 788 278 791
rect 214 751 217 758
rect 286 742 289 928
rect 294 872 297 908
rect 302 902 305 928
rect 310 902 313 948
rect 318 942 321 948
rect 334 932 337 938
rect 342 902 345 938
rect 358 932 361 938
rect 374 902 377 938
rect 398 932 401 958
rect 414 952 417 958
rect 414 938 422 941
rect 374 882 377 888
rect 386 868 390 871
rect 342 862 345 868
rect 358 862 361 868
rect 310 792 313 798
rect 302 762 305 768
rect 246 732 249 738
rect 214 672 217 728
rect 286 702 289 738
rect 246 692 249 698
rect 294 682 297 718
rect 270 672 273 678
rect 258 668 262 671
rect 258 658 262 661
rect 278 652 281 678
rect 302 672 305 758
rect 362 748 366 751
rect 334 742 337 748
rect 318 722 321 728
rect 334 672 337 678
rect 286 652 289 668
rect 298 658 302 661
rect 322 658 326 661
rect 210 568 214 571
rect 226 558 230 561
rect 198 552 201 558
rect 246 552 249 578
rect 246 542 249 548
rect 170 458 174 461
rect 182 452 185 458
rect 190 442 193 468
rect 198 372 201 538
rect 238 472 241 488
rect 278 472 281 528
rect 222 462 225 468
rect 226 448 230 451
rect 158 352 161 358
rect 182 352 185 358
rect 222 352 225 438
rect 118 348 126 351
rect 146 348 150 351
rect 6 292 9 328
rect 62 272 65 338
rect 62 262 65 268
rect 70 263 73 318
rect 102 292 105 328
rect 70 258 73 259
rect 62 152 65 258
rect 118 162 121 348
rect 190 342 193 348
rect 170 338 174 341
rect 162 328 166 331
rect 130 318 134 321
rect 202 318 206 321
rect 134 262 137 268
rect 166 263 169 318
rect 166 258 169 259
rect 102 152 105 158
rect 138 148 142 151
rect 54 132 57 148
rect 62 92 65 148
rect 110 142 113 148
rect 150 142 153 228
rect 206 152 209 268
rect 222 262 225 348
rect 254 332 257 468
rect 274 459 278 462
rect 286 362 289 648
rect 302 622 305 658
rect 322 648 326 651
rect 310 642 313 648
rect 330 638 334 641
rect 350 572 353 728
rect 366 682 369 738
rect 370 659 374 661
rect 366 658 374 659
rect 382 592 385 868
rect 406 862 409 868
rect 390 842 393 858
rect 398 852 401 858
rect 414 822 417 938
rect 422 922 425 928
rect 422 882 425 918
rect 430 902 433 948
rect 438 892 441 958
rect 454 952 457 958
rect 478 952 481 978
rect 494 952 497 968
rect 458 938 462 941
rect 474 938 486 941
rect 446 922 449 938
rect 498 888 502 891
rect 422 802 425 878
rect 438 872 441 878
rect 454 872 457 888
rect 454 862 457 868
rect 454 792 457 858
rect 510 821 513 938
rect 526 822 529 1058
rect 566 1042 569 1058
rect 558 962 561 1028
rect 582 1022 585 1058
rect 582 972 585 1018
rect 606 1012 609 1068
rect 578 958 585 961
rect 582 952 585 958
rect 554 948 558 951
rect 574 942 577 948
rect 586 938 590 941
rect 534 932 537 938
rect 598 922 601 938
rect 614 932 617 1068
rect 638 1062 641 1128
rect 646 1102 649 1158
rect 654 1122 657 1238
rect 678 1232 681 1248
rect 678 1152 681 1228
rect 686 1212 689 1248
rect 742 1242 745 1338
rect 758 1322 761 1328
rect 750 1301 753 1318
rect 766 1312 769 1338
rect 814 1322 817 1338
rect 750 1298 761 1301
rect 758 1252 761 1298
rect 782 1272 785 1308
rect 770 1258 774 1261
rect 782 1232 785 1268
rect 806 1262 809 1318
rect 822 1302 825 1318
rect 854 1282 857 1418
rect 838 1262 841 1278
rect 862 1272 865 1468
rect 950 1462 953 1488
rect 958 1462 961 1468
rect 998 1462 1001 1518
rect 1016 1503 1018 1507
rect 1022 1503 1025 1507
rect 1029 1503 1032 1507
rect 870 1432 873 1458
rect 894 1432 897 1448
rect 918 1372 921 1418
rect 1014 1372 1017 1468
rect 1046 1462 1049 1468
rect 1054 1462 1057 1668
rect 1070 1662 1073 1668
rect 1142 1662 1145 1668
rect 1158 1662 1161 1668
rect 1190 1662 1193 1718
rect 1214 1682 1217 1728
rect 1226 1718 1230 1721
rect 1254 1682 1257 1728
rect 1262 1692 1265 1698
rect 1242 1678 1246 1681
rect 1238 1662 1241 1678
rect 1114 1658 1118 1661
rect 1186 1658 1190 1661
rect 1062 1642 1065 1648
rect 1070 1632 1073 1648
rect 1086 1642 1089 1648
rect 1086 1562 1089 1568
rect 1066 1548 1070 1551
rect 1070 1512 1073 1538
rect 1094 1522 1097 1658
rect 1122 1648 1126 1651
rect 1126 1582 1129 1648
rect 1142 1572 1145 1658
rect 1206 1652 1209 1658
rect 1214 1652 1217 1658
rect 1246 1652 1249 1668
rect 1254 1662 1257 1668
rect 1258 1648 1262 1651
rect 1150 1622 1153 1648
rect 1206 1642 1209 1648
rect 1170 1638 1174 1641
rect 1166 1632 1169 1638
rect 1150 1572 1153 1618
rect 1122 1548 1126 1551
rect 1102 1532 1105 1538
rect 1110 1522 1113 1548
rect 1134 1532 1137 1538
rect 1070 1462 1073 1508
rect 1094 1462 1097 1518
rect 1118 1472 1121 1498
rect 1142 1471 1145 1568
rect 1158 1562 1161 1618
rect 1166 1562 1169 1578
rect 1150 1542 1153 1548
rect 1138 1468 1145 1471
rect 1042 1458 1046 1461
rect 1062 1452 1065 1458
rect 1118 1452 1121 1468
rect 1142 1461 1145 1468
rect 1142 1458 1150 1461
rect 1174 1452 1177 1568
rect 1190 1552 1193 1558
rect 1190 1522 1193 1548
rect 1182 1472 1185 1518
rect 1198 1512 1201 1538
rect 1206 1482 1209 1638
rect 1230 1612 1233 1618
rect 1246 1592 1249 1648
rect 1214 1562 1217 1588
rect 1214 1542 1217 1558
rect 1218 1538 1222 1541
rect 1234 1518 1238 1521
rect 1214 1482 1217 1518
rect 1026 1448 1030 1451
rect 1146 1448 1150 1451
rect 1174 1442 1177 1448
rect 1038 1402 1041 1438
rect 1070 1432 1073 1438
rect 1078 1402 1081 1438
rect 1094 1392 1097 1418
rect 886 1351 889 1358
rect 934 1342 937 1358
rect 1022 1352 1025 1358
rect 942 1342 945 1348
rect 870 1312 873 1338
rect 918 1302 921 1338
rect 870 1282 873 1298
rect 898 1288 902 1291
rect 882 1278 886 1281
rect 826 1248 830 1251
rect 846 1242 849 1268
rect 926 1262 929 1308
rect 858 1258 862 1261
rect 930 1258 937 1261
rect 946 1258 950 1261
rect 862 1242 865 1258
rect 670 1092 673 1098
rect 646 1082 649 1088
rect 666 1078 673 1081
rect 670 1072 673 1078
rect 678 1072 681 1118
rect 702 1112 705 1148
rect 718 1092 721 1098
rect 694 1072 697 1078
rect 622 992 625 998
rect 646 952 649 998
rect 654 972 657 1018
rect 670 992 673 1068
rect 702 1062 705 1088
rect 726 1081 729 1218
rect 750 1192 753 1218
rect 770 1148 774 1151
rect 726 1078 734 1081
rect 718 1062 721 1078
rect 726 1062 729 1068
rect 690 1058 694 1061
rect 658 948 662 951
rect 642 938 646 941
rect 614 912 617 928
rect 558 882 561 908
rect 590 872 593 888
rect 554 859 558 862
rect 606 862 609 868
rect 630 862 633 878
rect 638 872 641 888
rect 646 862 649 918
rect 662 892 665 898
rect 670 862 673 908
rect 678 892 681 1048
rect 694 992 697 1038
rect 718 1002 721 1058
rect 742 1031 745 1138
rect 766 1132 769 1148
rect 782 1082 785 1228
rect 790 1192 793 1228
rect 838 1201 841 1218
rect 838 1198 849 1201
rect 798 1142 801 1148
rect 750 1062 753 1068
rect 734 1028 745 1031
rect 734 1022 737 1028
rect 718 942 721 988
rect 734 952 737 1018
rect 742 982 745 1018
rect 758 952 761 1008
rect 766 962 769 968
rect 782 952 785 988
rect 790 972 793 1118
rect 822 1102 825 1118
rect 830 1092 833 1138
rect 838 1132 841 1188
rect 846 1141 849 1198
rect 862 1181 865 1218
rect 858 1178 865 1181
rect 862 1152 865 1158
rect 870 1152 873 1178
rect 918 1162 921 1168
rect 878 1152 881 1158
rect 862 1142 865 1148
rect 934 1142 937 1258
rect 958 1152 961 1348
rect 970 1338 974 1341
rect 982 1322 985 1328
rect 1016 1303 1018 1307
rect 1022 1303 1025 1307
rect 1029 1303 1032 1307
rect 990 1272 993 1288
rect 998 1268 1006 1271
rect 998 1262 1001 1268
rect 1006 1252 1009 1258
rect 966 1152 969 1158
rect 846 1138 854 1141
rect 798 1062 801 1078
rect 790 961 793 968
rect 790 958 798 961
rect 786 948 790 951
rect 742 942 745 948
rect 690 918 694 921
rect 718 892 721 938
rect 726 912 729 938
rect 734 872 737 918
rect 750 892 753 948
rect 786 938 790 941
rect 758 932 761 938
rect 742 882 745 888
rect 806 872 809 1008
rect 814 982 817 988
rect 830 962 833 968
rect 838 951 841 1128
rect 850 1088 854 1091
rect 854 1062 857 1068
rect 870 1062 873 1068
rect 878 1062 881 1088
rect 886 1082 889 1138
rect 894 1082 897 1138
rect 902 1092 905 1138
rect 942 1082 945 1088
rect 974 1082 977 1128
rect 898 1078 902 1081
rect 930 1068 934 1071
rect 894 1062 897 1068
rect 962 1058 966 1061
rect 906 1048 910 1051
rect 854 1042 857 1048
rect 834 948 841 951
rect 850 948 854 951
rect 862 942 865 968
rect 886 952 889 1018
rect 902 992 905 1038
rect 910 1032 913 1048
rect 918 1042 921 1058
rect 814 938 822 941
rect 754 868 758 871
rect 630 852 633 858
rect 610 848 614 851
rect 646 832 649 858
rect 510 818 521 821
rect 496 803 498 807
rect 502 803 505 807
rect 509 803 512 807
rect 422 772 425 778
rect 298 548 302 551
rect 330 488 334 491
rect 342 472 345 568
rect 398 562 401 768
rect 422 742 425 768
rect 442 758 446 761
rect 478 752 481 798
rect 502 762 505 788
rect 490 758 497 761
rect 506 758 510 761
rect 494 752 497 758
rect 466 748 470 751
rect 438 742 441 748
rect 478 742 481 748
rect 466 738 470 741
rect 478 732 481 738
rect 438 672 441 728
rect 462 692 465 698
rect 486 692 489 748
rect 510 742 513 748
rect 518 712 521 818
rect 534 782 537 788
rect 526 752 529 778
rect 550 762 553 768
rect 482 678 486 681
rect 498 678 502 681
rect 426 668 430 671
rect 474 668 478 671
rect 522 668 526 671
rect 510 662 513 668
rect 418 638 422 641
rect 414 592 417 628
rect 446 612 449 658
rect 462 652 465 658
rect 370 558 374 561
rect 378 548 382 551
rect 390 542 393 548
rect 398 542 401 558
rect 414 552 417 578
rect 430 562 433 588
rect 390 512 393 538
rect 318 372 321 378
rect 342 361 345 468
rect 350 462 353 478
rect 390 472 393 478
rect 370 468 374 471
rect 374 452 377 458
rect 406 422 409 538
rect 422 463 425 468
rect 422 458 425 459
rect 334 358 345 361
rect 274 348 278 351
rect 326 342 329 358
rect 334 352 337 358
rect 346 348 350 351
rect 230 262 233 278
rect 254 272 257 328
rect 286 292 289 308
rect 302 172 305 338
rect 334 322 337 348
rect 358 342 361 368
rect 374 362 377 368
rect 382 332 385 388
rect 430 371 433 558
rect 462 542 465 638
rect 470 582 473 658
rect 526 642 529 648
rect 496 603 498 607
rect 502 603 505 607
rect 509 603 512 607
rect 470 552 473 568
rect 446 462 449 538
rect 454 472 457 478
rect 510 472 513 558
rect 526 552 529 568
rect 534 542 537 738
rect 542 662 545 758
rect 582 752 585 818
rect 582 702 585 748
rect 590 742 593 748
rect 606 742 609 748
rect 614 742 617 778
rect 654 752 657 828
rect 662 752 665 818
rect 678 762 681 838
rect 694 752 697 858
rect 702 812 705 868
rect 798 862 801 868
rect 738 858 742 861
rect 770 858 774 861
rect 806 852 809 858
rect 714 848 718 851
rect 782 842 785 848
rect 726 832 729 838
rect 726 792 729 808
rect 814 792 817 938
rect 834 928 838 931
rect 822 872 825 898
rect 834 888 838 891
rect 830 852 833 868
rect 838 852 841 858
rect 830 832 833 848
rect 770 788 774 791
rect 706 758 710 761
rect 674 748 678 751
rect 622 742 625 748
rect 630 742 633 748
rect 710 742 713 748
rect 718 742 721 758
rect 806 752 809 788
rect 838 752 841 768
rect 730 748 734 751
rect 762 748 766 751
rect 786 748 790 751
rect 658 738 662 741
rect 682 738 686 741
rect 606 722 609 728
rect 586 688 590 691
rect 646 682 649 738
rect 682 728 686 731
rect 714 688 718 691
rect 550 672 553 678
rect 542 652 545 658
rect 566 652 569 658
rect 554 648 558 651
rect 574 582 577 668
rect 582 642 585 648
rect 562 568 566 571
rect 558 552 561 558
rect 438 392 441 428
rect 510 422 513 468
rect 518 462 521 488
rect 534 452 537 488
rect 496 403 498 407
rect 502 403 505 407
rect 509 403 512 407
rect 422 368 433 371
rect 398 352 401 358
rect 406 342 409 348
rect 422 332 425 368
rect 458 358 462 361
rect 430 342 433 358
rect 478 352 481 358
rect 438 342 441 348
rect 462 332 465 348
rect 390 322 393 328
rect 470 322 473 338
rect 486 332 489 338
rect 414 302 417 318
rect 510 302 513 348
rect 518 342 521 378
rect 310 252 313 288
rect 322 278 326 281
rect 342 272 345 288
rect 438 282 441 288
rect 358 272 361 278
rect 450 268 454 271
rect 330 258 334 261
rect 250 168 254 171
rect 290 158 294 161
rect 262 152 265 158
rect 194 148 198 151
rect 274 148 278 151
rect 302 142 305 168
rect 318 152 321 168
rect 326 142 329 258
rect 342 172 345 268
rect 382 252 385 258
rect 378 188 382 191
rect 398 162 401 268
rect 462 262 465 288
rect 494 272 497 278
rect 458 258 462 261
rect 478 252 481 268
rect 502 252 505 268
rect 482 248 486 251
rect 454 242 457 248
rect 496 203 498 207
rect 502 203 505 207
rect 509 203 512 207
rect 498 178 502 181
rect 342 152 345 158
rect 382 142 385 148
rect 98 138 102 141
rect 258 138 262 141
rect 314 138 318 141
rect 150 132 153 138
rect 358 132 361 138
rect 366 132 369 138
rect 398 132 401 158
rect 442 148 446 151
rect 518 142 521 168
rect 526 152 529 448
rect 542 441 545 468
rect 550 452 553 538
rect 566 492 569 528
rect 574 512 577 578
rect 582 562 585 568
rect 590 551 593 678
rect 598 612 601 668
rect 606 562 609 588
rect 582 548 593 551
rect 542 438 553 441
rect 534 392 537 438
rect 550 392 553 438
rect 566 432 569 448
rect 574 402 577 458
rect 582 392 585 548
rect 598 542 601 548
rect 590 492 593 508
rect 606 492 609 558
rect 614 472 617 668
rect 654 662 657 688
rect 698 678 702 681
rect 730 678 734 681
rect 706 668 710 671
rect 706 658 710 661
rect 734 652 737 678
rect 742 632 745 748
rect 750 742 753 748
rect 822 742 825 748
rect 786 738 790 741
rect 758 732 761 738
rect 798 732 801 738
rect 830 732 833 738
rect 790 692 793 698
rect 750 662 753 668
rect 758 662 761 688
rect 622 592 625 608
rect 630 572 633 578
rect 630 552 633 568
rect 622 542 625 548
rect 654 542 657 548
rect 634 538 638 541
rect 646 482 649 538
rect 662 532 665 618
rect 706 548 710 551
rect 750 542 753 658
rect 774 632 777 638
rect 790 602 793 648
rect 762 578 766 581
rect 766 558 774 561
rect 766 552 769 558
rect 798 552 801 558
rect 710 472 713 538
rect 766 532 769 538
rect 614 462 617 468
rect 710 462 713 468
rect 750 462 753 478
rect 774 472 777 548
rect 806 541 809 728
rect 838 721 841 738
rect 830 718 841 721
rect 814 652 817 658
rect 798 538 809 541
rect 814 542 817 578
rect 830 572 833 718
rect 846 692 849 928
rect 854 912 857 938
rect 870 902 873 948
rect 918 942 921 978
rect 934 962 937 988
rect 930 948 934 951
rect 906 938 913 941
rect 910 932 913 938
rect 898 928 902 931
rect 886 912 889 918
rect 898 888 902 891
rect 854 862 857 888
rect 934 882 937 918
rect 874 868 878 871
rect 922 868 926 871
rect 862 842 865 868
rect 862 762 865 778
rect 842 668 846 671
rect 854 661 857 718
rect 870 692 873 858
rect 910 842 913 858
rect 942 852 945 1018
rect 966 961 969 1018
rect 974 992 977 1048
rect 982 1042 985 1068
rect 998 1052 1001 1068
rect 958 958 969 961
rect 958 952 961 958
rect 966 942 969 948
rect 966 872 969 938
rect 942 822 945 848
rect 966 842 969 868
rect 918 792 921 818
rect 934 772 937 818
rect 878 731 881 758
rect 886 742 889 758
rect 894 742 897 748
rect 910 742 913 748
rect 902 731 905 738
rect 878 728 905 731
rect 882 718 886 721
rect 878 692 881 708
rect 870 672 873 678
rect 902 662 905 718
rect 918 662 921 768
rect 930 748 934 751
rect 934 692 937 738
rect 942 732 945 808
rect 958 772 961 818
rect 974 802 977 918
rect 982 882 985 1038
rect 990 952 993 978
rect 990 942 993 948
rect 990 862 993 868
rect 998 782 1001 938
rect 1006 882 1009 1248
rect 1022 1132 1025 1138
rect 1022 1122 1025 1128
rect 1016 1103 1018 1107
rect 1022 1103 1025 1107
rect 1029 1103 1032 1107
rect 1038 1062 1041 1378
rect 1054 1352 1057 1378
rect 1090 1348 1094 1351
rect 1046 1312 1049 1338
rect 1050 1268 1054 1271
rect 1050 1258 1054 1261
rect 1062 1252 1065 1348
rect 1102 1342 1105 1438
rect 1158 1402 1161 1438
rect 1182 1432 1185 1458
rect 1190 1442 1193 1478
rect 1218 1458 1222 1461
rect 1238 1452 1241 1508
rect 1246 1502 1249 1558
rect 1254 1492 1257 1518
rect 1206 1442 1209 1448
rect 1226 1438 1230 1441
rect 1246 1432 1249 1458
rect 1254 1452 1257 1488
rect 1270 1462 1273 1718
rect 1286 1672 1289 1718
rect 1406 1702 1409 1738
rect 1438 1682 1441 1728
rect 1342 1672 1345 1678
rect 1278 1462 1281 1578
rect 1286 1512 1289 1658
rect 1294 1562 1297 1668
rect 1454 1642 1457 1668
rect 1486 1662 1489 1738
rect 1322 1638 1326 1641
rect 1502 1622 1505 1648
rect 1398 1562 1401 1588
rect 1294 1462 1297 1558
rect 1334 1532 1337 1538
rect 1334 1492 1337 1508
rect 1350 1502 1353 1538
rect 1382 1532 1385 1548
rect 1470 1532 1473 1548
rect 1510 1542 1513 1728
rect 1558 1691 1561 1738
rect 1574 1732 1577 1738
rect 1614 1692 1617 1748
rect 1666 1738 1670 1741
rect 1734 1732 1737 1738
rect 1558 1688 1566 1691
rect 1542 1662 1545 1668
rect 1590 1662 1593 1668
rect 1528 1603 1530 1607
rect 1534 1603 1537 1607
rect 1541 1603 1544 1607
rect 1574 1562 1577 1588
rect 1582 1552 1585 1558
rect 1510 1532 1513 1538
rect 1434 1518 1438 1521
rect 1358 1482 1361 1508
rect 1406 1492 1409 1498
rect 1306 1478 1310 1481
rect 1370 1468 1374 1471
rect 1370 1458 1374 1461
rect 1270 1452 1273 1458
rect 1278 1452 1281 1458
rect 1258 1438 1262 1441
rect 1110 1352 1113 1378
rect 1134 1362 1137 1378
rect 1102 1322 1105 1338
rect 1074 1318 1078 1321
rect 1086 1272 1089 1278
rect 1094 1272 1097 1278
rect 1102 1272 1105 1278
rect 1074 1268 1078 1271
rect 1110 1262 1113 1348
rect 1126 1262 1129 1318
rect 1078 1252 1081 1258
rect 1062 1232 1065 1248
rect 1078 1192 1081 1248
rect 1102 1232 1105 1258
rect 1118 1222 1121 1258
rect 1134 1242 1137 1258
rect 1142 1192 1145 1348
rect 1150 1302 1153 1338
rect 1158 1312 1161 1318
rect 1150 1282 1153 1298
rect 1158 1282 1161 1288
rect 1166 1242 1169 1418
rect 1182 1412 1185 1418
rect 1230 1412 1233 1418
rect 1262 1372 1265 1418
rect 1190 1352 1193 1368
rect 1254 1362 1257 1368
rect 1218 1347 1222 1350
rect 1270 1342 1273 1428
rect 1278 1382 1281 1418
rect 1286 1392 1289 1438
rect 1294 1362 1297 1448
rect 1310 1412 1313 1418
rect 1318 1362 1321 1458
rect 1350 1442 1353 1458
rect 1382 1422 1385 1468
rect 1430 1451 1433 1488
rect 1462 1482 1465 1518
rect 1526 1492 1529 1538
rect 1598 1502 1601 1668
rect 1614 1642 1617 1658
rect 1646 1642 1649 1668
rect 1654 1642 1657 1718
rect 1670 1662 1673 1688
rect 1734 1682 1737 1728
rect 1670 1622 1673 1648
rect 1718 1602 1721 1668
rect 1630 1562 1633 1588
rect 1734 1582 1737 1678
rect 1774 1662 1777 1748
rect 1806 1692 1809 1738
rect 1822 1732 1825 1738
rect 1930 1728 1934 1731
rect 1902 1712 1905 1718
rect 1850 1688 1854 1691
rect 1902 1682 1905 1688
rect 1918 1681 1921 1718
rect 1942 1692 1945 1748
rect 1950 1732 1953 1738
rect 1958 1712 1961 1828
rect 2006 1762 2009 1768
rect 2046 1742 2049 1748
rect 2010 1728 2014 1731
rect 1966 1722 1969 1728
rect 1914 1678 1921 1681
rect 1878 1672 1881 1678
rect 1834 1668 1838 1671
rect 1914 1668 1918 1671
rect 1894 1662 1897 1668
rect 1870 1652 1873 1658
rect 1842 1648 1846 1651
rect 1798 1592 1801 1648
rect 1626 1548 1630 1551
rect 1678 1522 1681 1538
rect 1694 1532 1697 1538
rect 1734 1532 1737 1578
rect 1790 1552 1793 1558
rect 1782 1548 1790 1551
rect 1766 1518 1774 1521
rect 1546 1488 1550 1491
rect 1514 1478 1518 1481
rect 1462 1472 1465 1478
rect 1598 1472 1601 1498
rect 1610 1478 1614 1481
rect 1546 1468 1553 1471
rect 1438 1462 1441 1468
rect 1430 1448 1441 1451
rect 1414 1392 1417 1398
rect 1318 1352 1321 1358
rect 1342 1352 1345 1358
rect 1306 1348 1310 1351
rect 1362 1348 1366 1351
rect 1378 1348 1382 1351
rect 1174 1262 1177 1308
rect 1182 1292 1185 1298
rect 1238 1272 1241 1338
rect 1342 1332 1345 1338
rect 1258 1328 1262 1331
rect 1322 1328 1326 1331
rect 1350 1312 1353 1328
rect 1310 1262 1313 1278
rect 1234 1258 1238 1261
rect 1170 1228 1174 1231
rect 1054 1142 1057 1158
rect 1062 1142 1065 1158
rect 1078 1142 1081 1148
rect 1086 1142 1089 1188
rect 1190 1162 1193 1168
rect 1094 1152 1097 1158
rect 1046 1138 1054 1141
rect 1114 1138 1118 1141
rect 1178 1138 1182 1141
rect 1046 1072 1049 1138
rect 1022 1012 1025 1058
rect 1030 1052 1033 1058
rect 1022 952 1025 1008
rect 1016 903 1018 907
rect 1022 903 1025 907
rect 1029 903 1032 907
rect 1038 882 1041 1058
rect 1050 1038 1054 1041
rect 1078 952 1081 968
rect 1086 952 1089 1138
rect 1126 1122 1129 1138
rect 1134 1072 1137 1078
rect 1150 1062 1153 1118
rect 1198 1101 1201 1238
rect 1210 1158 1214 1161
rect 1206 1122 1209 1148
rect 1198 1098 1209 1101
rect 1206 1082 1209 1098
rect 1206 1072 1209 1078
rect 1214 1062 1217 1088
rect 1106 1058 1110 1061
rect 1134 952 1137 968
rect 1054 892 1057 948
rect 1054 872 1057 888
rect 1102 872 1105 948
rect 1142 942 1145 1028
rect 1150 982 1153 1058
rect 1170 1028 1174 1031
rect 1166 962 1169 978
rect 1154 948 1158 951
rect 1006 852 1009 858
rect 1030 852 1033 868
rect 1062 862 1065 868
rect 1042 858 1046 861
rect 1046 762 1049 858
rect 1102 852 1105 858
rect 1090 758 1094 761
rect 962 748 966 751
rect 974 742 977 758
rect 1118 752 1121 758
rect 978 738 982 741
rect 954 728 958 731
rect 990 682 993 688
rect 930 668 934 671
rect 986 668 990 671
rect 850 658 857 661
rect 838 542 841 648
rect 846 642 849 648
rect 862 642 865 658
rect 902 652 905 658
rect 934 652 937 658
rect 962 648 966 651
rect 850 638 857 641
rect 854 632 857 638
rect 846 552 849 568
rect 854 562 857 628
rect 878 622 881 648
rect 870 592 873 598
rect 594 358 598 361
rect 558 352 561 358
rect 614 352 617 378
rect 654 362 657 458
rect 694 422 697 428
rect 686 362 689 388
rect 634 358 638 361
rect 646 352 649 358
rect 670 352 673 358
rect 658 348 662 351
rect 686 342 689 358
rect 658 338 662 341
rect 694 341 697 418
rect 750 412 753 438
rect 734 352 737 398
rect 750 392 753 408
rect 798 392 801 538
rect 814 528 822 531
rect 806 462 809 468
rect 806 362 809 368
rect 694 338 702 341
rect 534 332 537 338
rect 582 332 585 338
rect 542 312 545 328
rect 550 272 553 298
rect 558 262 561 268
rect 546 258 550 261
rect 566 182 569 328
rect 574 252 577 328
rect 590 292 593 308
rect 614 302 617 338
rect 606 298 614 301
rect 590 192 593 258
rect 598 232 601 268
rect 606 262 609 298
rect 614 272 617 278
rect 622 261 625 338
rect 630 272 633 278
rect 670 272 673 298
rect 694 292 697 318
rect 718 302 721 318
rect 750 292 753 358
rect 814 352 817 528
rect 830 522 833 528
rect 838 512 841 518
rect 846 512 849 548
rect 870 532 873 548
rect 886 542 889 608
rect 914 558 918 561
rect 894 552 897 558
rect 926 551 929 558
rect 918 548 929 551
rect 966 551 969 558
rect 918 542 921 548
rect 878 532 881 538
rect 934 532 937 538
rect 822 472 825 478
rect 822 452 825 458
rect 822 412 825 448
rect 830 402 833 478
rect 774 342 777 348
rect 798 332 801 348
rect 658 268 662 271
rect 722 268 726 271
rect 622 258 630 261
rect 622 232 625 258
rect 634 248 638 251
rect 654 242 657 248
rect 550 162 553 168
rect 534 142 537 148
rect 566 142 569 178
rect 606 151 609 228
rect 662 222 665 258
rect 622 192 625 218
rect 678 192 681 258
rect 694 252 697 268
rect 730 258 734 261
rect 742 252 745 258
rect 722 248 726 251
rect 602 148 609 151
rect 614 142 617 148
rect 114 128 118 131
rect 390 122 393 128
rect 246 82 249 98
rect 10 68 14 71
rect 74 68 78 71
rect 142 62 145 68
rect 158 62 161 68
rect 262 62 265 108
rect 286 72 289 108
rect 270 62 273 68
rect 310 62 313 68
rect 334 62 337 118
rect 390 92 393 118
rect 186 58 190 61
rect 290 58 294 61
rect 398 52 401 118
rect 414 101 417 128
rect 414 98 425 101
rect 414 62 417 88
rect 422 72 425 98
rect 430 92 433 138
rect 438 62 441 138
rect 574 122 577 128
rect 614 82 617 128
rect 598 72 601 78
rect 654 62 657 68
rect 678 62 681 168
rect 686 151 689 228
rect 694 192 697 248
rect 702 242 705 248
rect 726 152 729 168
rect 758 161 761 328
rect 782 322 785 328
rect 822 322 825 348
rect 838 342 841 508
rect 870 492 873 498
rect 878 482 881 488
rect 846 462 849 468
rect 886 462 889 508
rect 902 492 905 528
rect 910 482 913 488
rect 918 472 921 508
rect 946 488 950 491
rect 958 472 961 498
rect 846 352 849 388
rect 854 372 857 458
rect 862 452 865 458
rect 894 432 897 468
rect 926 462 929 468
rect 950 452 953 468
rect 974 462 977 468
rect 982 462 985 598
rect 998 552 1001 738
rect 1022 732 1025 748
rect 1126 742 1129 938
rect 1158 932 1161 938
rect 1158 882 1161 888
rect 1166 871 1169 958
rect 1182 951 1185 968
rect 1222 962 1225 1238
rect 1230 1192 1233 1218
rect 1238 1152 1241 1198
rect 1294 1172 1297 1178
rect 1298 1148 1302 1151
rect 1238 1102 1241 1138
rect 1246 1112 1249 1148
rect 1310 1142 1313 1248
rect 1350 1242 1353 1248
rect 1326 1162 1329 1168
rect 1298 1138 1302 1141
rect 1322 1138 1326 1141
rect 1254 992 1257 1138
rect 1310 1132 1313 1138
rect 1266 1128 1270 1131
rect 1338 1118 1342 1121
rect 1270 1092 1273 1108
rect 1238 982 1241 988
rect 1194 958 1198 961
rect 1222 952 1225 958
rect 1262 952 1265 1008
rect 1278 1002 1281 1098
rect 1314 1088 1318 1091
rect 1322 1068 1326 1071
rect 1294 1062 1297 1068
rect 1278 992 1281 998
rect 1182 948 1193 951
rect 1174 942 1177 948
rect 1190 942 1193 948
rect 1226 938 1230 941
rect 1254 922 1257 948
rect 1254 902 1257 918
rect 1270 872 1273 938
rect 1302 932 1305 938
rect 1318 902 1321 1068
rect 1342 1062 1345 1078
rect 1358 1072 1361 1348
rect 1366 1342 1369 1348
rect 1386 1338 1390 1341
rect 1398 1302 1401 1348
rect 1370 1288 1374 1291
rect 1390 1272 1393 1278
rect 1378 1268 1382 1271
rect 1406 1262 1409 1378
rect 1422 1352 1425 1438
rect 1438 1352 1441 1448
rect 1466 1448 1470 1451
rect 1454 1432 1457 1448
rect 1486 1442 1489 1458
rect 1494 1422 1497 1468
rect 1446 1372 1449 1418
rect 1454 1392 1457 1418
rect 1528 1403 1530 1407
rect 1534 1403 1537 1407
rect 1541 1403 1544 1407
rect 1550 1392 1553 1468
rect 1558 1412 1561 1468
rect 1574 1452 1577 1458
rect 1590 1452 1593 1458
rect 1614 1392 1617 1418
rect 1486 1362 1489 1388
rect 1614 1362 1617 1378
rect 1490 1358 1494 1361
rect 1614 1352 1617 1358
rect 1426 1348 1430 1351
rect 1462 1342 1465 1348
rect 1526 1342 1529 1348
rect 1462 1312 1465 1338
rect 1566 1322 1569 1348
rect 1630 1332 1633 1498
rect 1698 1488 1702 1491
rect 1638 1442 1641 1448
rect 1646 1372 1649 1468
rect 1670 1422 1673 1448
rect 1662 1352 1665 1358
rect 1642 1348 1646 1351
rect 1654 1332 1657 1348
rect 1614 1321 1617 1328
rect 1638 1321 1641 1328
rect 1614 1318 1641 1321
rect 1450 1288 1454 1291
rect 1422 1272 1425 1288
rect 1542 1282 1545 1288
rect 1578 1268 1582 1271
rect 1510 1263 1513 1268
rect 1386 1258 1390 1261
rect 1598 1262 1601 1268
rect 1606 1262 1609 1298
rect 1618 1278 1622 1281
rect 1646 1272 1649 1278
rect 1618 1268 1622 1271
rect 1578 1258 1582 1261
rect 1406 1252 1409 1258
rect 1478 1252 1481 1258
rect 1382 1152 1385 1158
rect 1422 1132 1425 1248
rect 1438 1162 1441 1218
rect 1446 1202 1449 1218
rect 1470 1160 1473 1179
rect 1438 1142 1441 1148
rect 1378 1078 1382 1081
rect 1478 1072 1481 1248
rect 1598 1212 1601 1258
rect 1528 1203 1530 1207
rect 1534 1203 1537 1207
rect 1541 1203 1544 1207
rect 1494 1152 1497 1178
rect 1622 1172 1625 1258
rect 1630 1232 1633 1268
rect 1662 1262 1665 1348
rect 1678 1342 1681 1478
rect 1686 1472 1689 1478
rect 1710 1472 1713 1488
rect 1734 1472 1737 1488
rect 1742 1482 1745 1488
rect 1710 1422 1713 1458
rect 1718 1452 1721 1468
rect 1766 1462 1769 1518
rect 1774 1512 1777 1518
rect 1782 1502 1785 1548
rect 1806 1532 1809 1548
rect 1802 1528 1806 1531
rect 1774 1472 1777 1478
rect 1726 1412 1729 1418
rect 1702 1362 1705 1378
rect 1718 1352 1721 1408
rect 1734 1401 1737 1448
rect 1730 1398 1737 1401
rect 1726 1362 1729 1378
rect 1750 1372 1753 1428
rect 1766 1412 1769 1458
rect 1782 1431 1785 1498
rect 1790 1462 1793 1528
rect 1814 1492 1817 1618
rect 1846 1562 1849 1568
rect 1834 1538 1838 1541
rect 1822 1491 1825 1518
rect 1830 1502 1833 1528
rect 1838 1492 1841 1518
rect 1846 1512 1849 1548
rect 1870 1532 1873 1558
rect 1886 1552 1889 1658
rect 1966 1642 1969 1668
rect 1974 1652 1977 1668
rect 1982 1662 1985 1678
rect 1994 1658 1998 1661
rect 2006 1652 2009 1708
rect 2014 1652 2017 1658
rect 1914 1558 1918 1561
rect 1902 1552 1905 1558
rect 1934 1552 1937 1558
rect 1894 1542 1897 1548
rect 1958 1542 1961 1578
rect 1874 1528 1878 1531
rect 1886 1531 1889 1538
rect 1886 1528 1897 1531
rect 1822 1488 1833 1491
rect 1830 1482 1833 1488
rect 1878 1482 1881 1518
rect 1894 1492 1897 1528
rect 1918 1502 1921 1518
rect 1942 1512 1945 1538
rect 1966 1492 1969 1508
rect 1910 1482 1913 1488
rect 1954 1478 1958 1481
rect 1790 1452 1793 1458
rect 1774 1428 1785 1431
rect 1758 1382 1761 1388
rect 1738 1348 1742 1351
rect 1674 1318 1678 1321
rect 1686 1302 1689 1348
rect 1750 1342 1753 1368
rect 1694 1282 1697 1288
rect 1690 1268 1694 1271
rect 1674 1258 1678 1261
rect 1630 1192 1633 1208
rect 1518 1162 1521 1168
rect 1570 1148 1574 1151
rect 1510 1111 1513 1148
rect 1598 1142 1601 1158
rect 1606 1142 1609 1148
rect 1622 1142 1625 1168
rect 1638 1162 1641 1258
rect 1650 1248 1654 1251
rect 1654 1192 1657 1238
rect 1702 1192 1705 1318
rect 1718 1312 1721 1338
rect 1766 1322 1769 1368
rect 1774 1352 1777 1428
rect 1782 1372 1785 1418
rect 1786 1358 1790 1361
rect 1798 1352 1801 1458
rect 1806 1442 1809 1448
rect 1806 1352 1809 1358
rect 1786 1348 1790 1351
rect 1786 1338 1790 1341
rect 1802 1338 1806 1341
rect 1814 1332 1817 1478
rect 1822 1472 1825 1478
rect 1846 1472 1849 1478
rect 1882 1468 1886 1471
rect 1822 1452 1825 1458
rect 1830 1402 1833 1468
rect 1866 1458 1870 1461
rect 1882 1458 1886 1461
rect 1846 1362 1849 1368
rect 1854 1352 1857 1458
rect 1866 1438 1870 1441
rect 1910 1432 1913 1478
rect 1942 1462 1945 1468
rect 1974 1462 1977 1468
rect 1926 1422 1929 1458
rect 1934 1442 1937 1448
rect 1946 1438 1950 1441
rect 1970 1438 1974 1441
rect 1910 1392 1913 1418
rect 1926 1392 1929 1398
rect 1934 1362 1937 1368
rect 1950 1362 1953 1428
rect 1958 1362 1961 1418
rect 1982 1362 1985 1548
rect 1998 1492 2001 1648
rect 2006 1532 2009 1648
rect 2022 1642 2025 1728
rect 2038 1682 2041 1688
rect 2046 1672 2049 1678
rect 2006 1511 2009 1528
rect 2006 1508 2017 1511
rect 1990 1432 1993 1448
rect 1998 1382 2001 1418
rect 1898 1358 1902 1361
rect 1834 1348 1838 1351
rect 1862 1342 1865 1348
rect 1838 1332 1841 1338
rect 1862 1322 1865 1338
rect 1710 1282 1713 1308
rect 1770 1288 1774 1291
rect 1798 1282 1801 1318
rect 1726 1262 1729 1268
rect 1734 1262 1737 1268
rect 1742 1262 1745 1278
rect 1742 1252 1745 1258
rect 1774 1252 1777 1278
rect 1714 1248 1718 1251
rect 1790 1242 1793 1268
rect 1798 1252 1801 1278
rect 1814 1272 1817 1288
rect 1838 1282 1841 1288
rect 1870 1272 1873 1298
rect 1878 1292 1881 1358
rect 1942 1342 1945 1348
rect 1922 1338 1926 1341
rect 1874 1268 1878 1271
rect 1886 1271 1889 1308
rect 1894 1302 1897 1338
rect 1950 1302 1953 1358
rect 1974 1342 1977 1358
rect 2006 1352 2009 1508
rect 2014 1470 2017 1508
rect 2022 1482 2025 1638
rect 2022 1472 2025 1478
rect 2014 1392 2017 1438
rect 2030 1371 2033 1418
rect 2038 1382 2041 1518
rect 2046 1462 2049 1668
rect 2030 1368 2038 1371
rect 1986 1348 1990 1351
rect 2046 1342 2049 1458
rect 1962 1338 1966 1341
rect 1986 1338 1990 1341
rect 2006 1332 2010 1335
rect 1958 1322 1961 1328
rect 1990 1292 1993 1298
rect 1902 1272 1905 1288
rect 1998 1282 2001 1298
rect 2030 1292 2033 1298
rect 2026 1278 2030 1281
rect 1886 1268 1894 1271
rect 1822 1252 1825 1258
rect 1854 1252 1857 1268
rect 1934 1262 1937 1278
rect 2014 1272 2017 1278
rect 1958 1262 1961 1268
rect 1938 1258 1942 1261
rect 1854 1242 1857 1248
rect 1670 1162 1673 1178
rect 1642 1158 1646 1161
rect 1630 1152 1633 1158
rect 1646 1142 1649 1148
rect 1570 1138 1574 1141
rect 1654 1132 1657 1148
rect 1502 1108 1513 1111
rect 1518 1128 1526 1131
rect 1370 1068 1374 1071
rect 1454 1062 1457 1068
rect 1370 1058 1374 1061
rect 1326 1022 1329 1058
rect 1334 1052 1337 1058
rect 1326 932 1329 948
rect 1166 868 1174 871
rect 1142 862 1145 868
rect 1222 862 1225 868
rect 1254 863 1257 868
rect 1186 858 1190 861
rect 1286 862 1289 878
rect 1302 862 1305 898
rect 1334 872 1337 898
rect 1314 868 1318 871
rect 1342 862 1345 918
rect 1350 892 1353 1048
rect 1366 1022 1369 1058
rect 1398 952 1401 1038
rect 1502 992 1505 1108
rect 1386 948 1390 951
rect 1418 948 1422 951
rect 1398 942 1401 948
rect 1382 922 1385 938
rect 1406 922 1409 928
rect 1374 892 1377 908
rect 1166 852 1169 858
rect 1190 842 1193 858
rect 1158 792 1161 828
rect 1146 788 1150 791
rect 1158 762 1161 788
rect 1074 738 1078 741
rect 1016 703 1018 707
rect 1022 703 1025 707
rect 1029 703 1032 707
rect 1014 582 1017 658
rect 1022 652 1025 658
rect 1030 572 1033 668
rect 1046 652 1049 738
rect 1134 732 1137 758
rect 1162 748 1166 751
rect 1150 732 1153 748
rect 1182 742 1185 778
rect 1194 768 1198 771
rect 1222 752 1225 858
rect 1302 752 1305 858
rect 1334 832 1337 858
rect 1250 747 1254 750
rect 1098 728 1102 731
rect 1062 672 1065 698
rect 1158 692 1161 728
rect 1182 682 1185 688
rect 1194 678 1198 681
rect 1230 672 1233 678
rect 1178 668 1190 671
rect 1106 658 1110 661
rect 1038 632 1041 648
rect 962 458 966 461
rect 938 448 942 451
rect 982 442 985 458
rect 894 392 897 398
rect 766 262 769 268
rect 774 262 777 298
rect 750 158 761 161
rect 774 162 777 238
rect 782 222 785 268
rect 798 252 801 268
rect 798 192 801 208
rect 722 138 726 141
rect 686 82 689 108
rect 702 82 705 138
rect 742 132 745 158
rect 750 142 753 158
rect 794 148 798 151
rect 686 72 689 78
rect 702 72 705 78
rect 742 62 745 118
rect 758 102 761 148
rect 790 92 793 128
rect 782 82 785 88
rect 806 82 809 318
rect 830 302 833 338
rect 834 298 841 301
rect 822 262 825 288
rect 830 272 833 278
rect 838 272 841 298
rect 846 272 849 348
rect 854 282 857 368
rect 870 362 873 388
rect 990 352 993 368
rect 934 342 937 348
rect 974 342 977 348
rect 866 338 870 341
rect 990 332 993 348
rect 998 342 1001 548
rect 1038 532 1041 628
rect 1030 522 1033 528
rect 1016 503 1018 507
rect 1022 503 1025 507
rect 1029 503 1032 507
rect 1038 472 1041 528
rect 1046 492 1049 558
rect 1054 522 1057 658
rect 1126 652 1129 658
rect 1070 592 1073 618
rect 1102 542 1105 558
rect 1118 552 1121 558
rect 1138 548 1142 551
rect 1150 542 1153 608
rect 1166 582 1169 658
rect 1246 652 1249 738
rect 1286 732 1289 738
rect 1294 682 1297 718
rect 1302 671 1305 748
rect 1310 732 1313 768
rect 1350 762 1353 888
rect 1422 882 1425 948
rect 1446 942 1449 988
rect 1454 942 1457 948
rect 1470 942 1473 958
rect 1438 932 1441 938
rect 1478 932 1481 948
rect 1486 942 1489 988
rect 1518 982 1521 1128
rect 1542 1032 1545 1128
rect 1558 1122 1561 1128
rect 1582 1122 1585 1128
rect 1590 1122 1593 1128
rect 1558 1062 1561 1098
rect 1622 1092 1625 1098
rect 1598 1082 1601 1088
rect 1638 1072 1641 1118
rect 1650 1078 1654 1081
rect 1610 1068 1614 1071
rect 1638 1062 1641 1068
rect 1662 1062 1665 1158
rect 1658 1058 1662 1061
rect 1606 1032 1609 1058
rect 1528 1003 1530 1007
rect 1534 1003 1537 1007
rect 1541 1003 1544 1007
rect 1510 942 1513 948
rect 1498 938 1502 941
rect 1518 941 1521 978
rect 1614 952 1617 968
rect 1634 958 1638 961
rect 1518 938 1526 941
rect 1470 902 1473 918
rect 1358 762 1361 818
rect 1326 752 1329 758
rect 1350 742 1353 758
rect 1346 728 1350 731
rect 1346 678 1350 681
rect 1326 672 1329 678
rect 1302 668 1310 671
rect 1262 663 1265 668
rect 1262 658 1265 659
rect 1190 562 1193 568
rect 1162 548 1166 551
rect 1238 542 1241 548
rect 1246 542 1249 648
rect 1278 622 1281 668
rect 1294 552 1297 668
rect 1358 662 1361 748
rect 1366 742 1369 878
rect 1486 871 1489 938
rect 1526 932 1529 938
rect 1506 928 1510 931
rect 1546 928 1550 931
rect 1502 892 1505 908
rect 1486 868 1494 871
rect 1438 863 1441 868
rect 1454 862 1457 868
rect 1502 862 1505 888
rect 1518 862 1521 888
rect 1566 882 1569 948
rect 1574 892 1577 938
rect 1606 932 1609 938
rect 1594 928 1598 931
rect 1614 922 1617 938
rect 1638 902 1641 958
rect 1662 952 1665 958
rect 1670 952 1673 1158
rect 1694 1152 1697 1168
rect 1710 1160 1713 1179
rect 1742 1142 1745 1238
rect 1758 1162 1761 1218
rect 1758 1132 1761 1138
rect 1730 1088 1734 1091
rect 1678 1082 1681 1088
rect 1710 1082 1713 1088
rect 1690 1078 1694 1081
rect 1762 1078 1766 1081
rect 1710 1062 1713 1078
rect 1750 1072 1753 1078
rect 1694 1002 1697 1058
rect 1678 962 1681 978
rect 1666 938 1670 941
rect 1678 932 1681 958
rect 1694 952 1697 958
rect 1702 942 1705 1058
rect 1726 1052 1729 1058
rect 1806 1052 1809 1218
rect 1886 1212 1889 1218
rect 1910 1212 1913 1218
rect 1838 1182 1841 1188
rect 1886 1142 1889 1148
rect 1910 1142 1913 1148
rect 1854 1102 1857 1118
rect 1838 1052 1841 1059
rect 1730 1048 1737 1051
rect 1718 962 1721 968
rect 1722 948 1729 951
rect 1558 878 1566 881
rect 1490 858 1494 861
rect 1514 858 1518 861
rect 1474 848 1478 851
rect 1374 752 1377 768
rect 1398 762 1401 768
rect 1414 742 1417 768
rect 1446 742 1449 747
rect 1366 722 1369 738
rect 1430 732 1433 738
rect 1394 728 1398 731
rect 1366 672 1369 718
rect 1398 692 1401 698
rect 1406 682 1409 688
rect 1374 662 1377 668
rect 1306 658 1310 661
rect 1318 562 1321 648
rect 1302 552 1305 558
rect 1318 542 1321 558
rect 1162 538 1166 541
rect 1290 538 1294 541
rect 1078 532 1081 538
rect 1126 522 1129 528
rect 1078 492 1081 498
rect 1086 482 1089 498
rect 1102 492 1105 518
rect 1094 482 1097 488
rect 1006 372 1009 468
rect 1030 452 1033 458
rect 1038 352 1041 438
rect 1046 392 1049 468
rect 1054 462 1057 478
rect 1110 472 1113 498
rect 1074 468 1078 471
rect 1122 468 1126 471
rect 1142 462 1145 488
rect 1150 472 1153 508
rect 1158 462 1161 538
rect 1178 528 1182 531
rect 1166 492 1169 528
rect 1174 512 1177 518
rect 1174 482 1177 498
rect 1222 462 1225 508
rect 1246 482 1249 538
rect 1066 458 1070 461
rect 1122 458 1126 461
rect 1054 432 1057 458
rect 1054 342 1057 348
rect 1006 322 1009 328
rect 1062 322 1065 338
rect 866 288 881 291
rect 878 282 881 288
rect 814 232 817 258
rect 814 152 817 198
rect 830 192 833 258
rect 862 252 865 268
rect 870 262 873 278
rect 950 272 953 278
rect 914 268 918 271
rect 938 268 942 271
rect 898 258 902 261
rect 930 258 934 261
rect 878 252 881 258
rect 858 158 862 161
rect 818 138 822 141
rect 806 72 809 78
rect 822 72 825 128
rect 838 102 841 138
rect 846 62 849 68
rect 862 62 865 118
rect 870 62 873 218
rect 878 152 881 158
rect 886 142 889 258
rect 902 252 905 258
rect 942 222 945 248
rect 894 212 897 218
rect 942 152 945 208
rect 958 192 961 258
rect 966 251 969 268
rect 974 262 977 268
rect 982 262 985 268
rect 990 262 993 318
rect 1016 303 1018 307
rect 1022 303 1025 307
rect 1029 303 1032 307
rect 1010 258 1014 261
rect 966 248 974 251
rect 990 192 993 258
rect 1006 212 1009 218
rect 998 142 1001 148
rect 878 138 886 141
rect 878 92 881 138
rect 982 132 985 138
rect 1006 132 1009 168
rect 1022 152 1025 178
rect 994 128 998 131
rect 910 92 913 98
rect 918 72 921 128
rect 1016 103 1018 107
rect 1022 103 1025 107
rect 1029 103 1032 107
rect 1038 92 1041 318
rect 1054 292 1057 318
rect 1046 272 1049 278
rect 1062 232 1065 268
rect 1070 262 1073 458
rect 1262 452 1265 468
rect 1278 462 1281 468
rect 1130 448 1134 451
rect 1090 368 1094 371
rect 1110 352 1113 398
rect 1118 352 1121 368
rect 1078 292 1081 348
rect 1102 342 1105 348
rect 1118 312 1121 348
rect 1130 338 1134 341
rect 1142 332 1145 448
rect 1278 442 1281 448
rect 1206 352 1209 368
rect 1154 338 1158 341
rect 1046 192 1049 228
rect 1026 88 1030 91
rect 1078 82 1081 288
rect 1118 272 1121 278
rect 1126 272 1129 318
rect 1134 272 1137 318
rect 1158 272 1161 328
rect 1190 272 1193 298
rect 1094 262 1097 268
rect 1126 252 1129 258
rect 1134 252 1137 258
rect 1102 152 1105 218
rect 1150 172 1153 258
rect 1158 212 1161 268
rect 1166 252 1169 268
rect 1214 262 1217 278
rect 1222 272 1225 428
rect 1246 342 1249 398
rect 1286 392 1289 538
rect 1294 462 1297 518
rect 1326 512 1329 658
rect 1338 648 1342 651
rect 1334 542 1337 548
rect 1350 542 1353 618
rect 1366 592 1369 658
rect 1374 652 1377 658
rect 1366 551 1369 558
rect 1334 482 1337 528
rect 1346 488 1350 491
rect 1302 462 1305 468
rect 1334 462 1337 478
rect 1382 462 1385 658
rect 1390 542 1393 668
rect 1414 662 1417 698
rect 1450 678 1454 681
rect 1446 662 1449 668
rect 1462 662 1465 678
rect 1470 672 1473 838
rect 1534 832 1537 858
rect 1486 792 1489 818
rect 1528 803 1530 807
rect 1534 803 1537 807
rect 1541 803 1544 807
rect 1506 768 1510 771
rect 1478 682 1481 758
rect 1494 692 1497 758
rect 1534 752 1537 788
rect 1546 738 1550 741
rect 1558 732 1561 878
rect 1582 872 1585 898
rect 1646 892 1649 918
rect 1590 872 1593 888
rect 1566 862 1569 868
rect 1646 862 1649 868
rect 1590 852 1593 858
rect 1566 732 1569 768
rect 1578 758 1582 761
rect 1610 758 1614 761
rect 1590 752 1593 758
rect 1598 742 1601 748
rect 1630 742 1633 808
rect 1578 738 1582 741
rect 1546 728 1550 731
rect 1478 672 1481 678
rect 1502 672 1505 678
rect 1534 672 1537 678
rect 1510 662 1513 668
rect 1518 662 1521 668
rect 1414 602 1417 658
rect 1478 652 1481 658
rect 1542 652 1545 688
rect 1606 682 1609 738
rect 1614 692 1617 718
rect 1630 682 1633 738
rect 1470 648 1478 651
rect 1470 592 1473 648
rect 1528 603 1530 607
rect 1534 603 1537 607
rect 1541 603 1544 607
rect 1506 548 1510 551
rect 1534 551 1537 588
rect 1398 472 1401 548
rect 1418 538 1422 541
rect 1438 532 1441 548
rect 1566 542 1569 668
rect 1582 663 1585 668
rect 1582 658 1585 659
rect 1590 552 1593 558
rect 1590 522 1593 548
rect 1454 492 1457 518
rect 1438 482 1441 488
rect 1498 478 1502 481
rect 1478 472 1481 478
rect 1518 472 1521 488
rect 1558 472 1561 478
rect 1598 472 1601 508
rect 1282 348 1286 351
rect 1302 342 1305 348
rect 1250 268 1254 271
rect 1262 271 1265 328
rect 1278 292 1281 338
rect 1298 318 1302 321
rect 1318 272 1321 418
rect 1398 402 1401 468
rect 1406 463 1409 468
rect 1454 462 1457 468
rect 1462 462 1465 468
rect 1326 352 1329 388
rect 1398 372 1401 398
rect 1370 368 1374 371
rect 1350 352 1353 368
rect 1358 352 1361 358
rect 1334 342 1337 348
rect 1422 342 1425 348
rect 1262 268 1270 271
rect 1274 268 1278 271
rect 1330 268 1334 271
rect 1318 262 1321 268
rect 1366 262 1369 318
rect 1422 282 1425 308
rect 1430 292 1433 328
rect 1446 282 1449 288
rect 1462 272 1465 338
rect 1478 272 1481 468
rect 1486 462 1489 468
rect 1598 462 1601 468
rect 1566 458 1574 461
rect 1490 448 1494 451
rect 1510 442 1513 458
rect 1558 452 1561 458
rect 1486 392 1489 428
rect 1528 403 1530 407
rect 1534 403 1537 407
rect 1541 403 1544 407
rect 1550 391 1553 418
rect 1546 388 1553 391
rect 1406 262 1409 268
rect 1202 258 1206 261
rect 1242 258 1246 261
rect 1266 258 1270 261
rect 1442 258 1446 261
rect 1190 232 1193 258
rect 1202 248 1206 251
rect 1250 248 1254 251
rect 1182 222 1185 228
rect 1294 212 1297 248
rect 1302 192 1305 238
rect 1154 158 1158 161
rect 1158 152 1161 158
rect 1174 152 1177 158
rect 1186 148 1190 151
rect 1222 151 1225 158
rect 1186 138 1190 141
rect 1102 122 1105 138
rect 1142 132 1145 138
rect 1206 122 1209 138
rect 1254 132 1257 138
rect 1102 72 1105 118
rect 1310 92 1313 258
rect 1366 152 1369 158
rect 1358 142 1361 148
rect 1374 92 1377 148
rect 1226 88 1230 91
rect 1330 88 1334 91
rect 1118 72 1121 88
rect 1190 82 1193 88
rect 1166 72 1169 78
rect 1214 72 1217 78
rect 1310 72 1313 78
rect 1374 72 1377 78
rect 942 62 945 68
rect 1054 62 1057 68
rect 1086 63 1089 68
rect 466 58 470 61
rect 578 58 582 61
rect 962 58 966 61
rect 1134 62 1137 68
rect 1166 62 1169 68
rect 1174 62 1177 68
rect 1390 62 1393 118
rect 1406 82 1409 258
rect 1462 242 1465 268
rect 1510 263 1513 298
rect 1542 262 1545 388
rect 1558 362 1561 448
rect 1566 442 1569 458
rect 1566 392 1569 438
rect 1590 382 1593 418
rect 1606 392 1609 678
rect 1638 652 1641 728
rect 1646 641 1649 858
rect 1654 762 1657 878
rect 1666 858 1670 861
rect 1678 782 1681 918
rect 1710 872 1713 938
rect 1710 862 1713 868
rect 1718 862 1721 918
rect 1714 848 1718 851
rect 1726 842 1729 948
rect 1734 932 1737 1048
rect 1822 992 1825 1038
rect 1802 958 1806 961
rect 1822 952 1825 988
rect 1854 972 1857 1068
rect 1870 1062 1873 1068
rect 1918 1062 1921 1258
rect 1974 1151 1977 1268
rect 1982 1242 1985 1268
rect 2002 1258 2006 1261
rect 1982 1122 1985 1238
rect 2038 1192 2041 1268
rect 2046 1242 2049 1258
rect 1926 1062 1929 1078
rect 1966 1072 1969 1108
rect 1990 1092 1993 1148
rect 2014 1072 2017 1098
rect 1970 1068 1974 1071
rect 1906 1058 1910 1061
rect 1954 1058 1958 1061
rect 1878 1042 1881 1058
rect 1902 1032 1905 1058
rect 1894 952 1897 1018
rect 1754 938 1758 941
rect 1738 928 1742 931
rect 1742 852 1745 898
rect 1766 892 1769 948
rect 1774 912 1777 948
rect 1782 922 1785 948
rect 1758 872 1761 888
rect 1782 862 1785 898
rect 1794 888 1798 891
rect 1790 872 1793 878
rect 1770 858 1774 861
rect 1710 792 1713 838
rect 1654 752 1657 758
rect 1678 742 1681 758
rect 1686 722 1689 748
rect 1694 732 1697 748
rect 1726 732 1729 768
rect 1734 752 1737 848
rect 1758 752 1761 768
rect 1806 752 1809 948
rect 1894 872 1897 938
rect 1902 862 1905 1008
rect 1910 862 1913 868
rect 1850 858 1854 861
rect 1830 772 1833 858
rect 1814 762 1817 768
rect 1770 748 1774 751
rect 1738 738 1742 741
rect 1758 732 1761 748
rect 1798 742 1801 748
rect 1786 738 1790 741
rect 1654 662 1657 668
rect 1662 662 1665 668
rect 1646 638 1654 641
rect 1630 492 1633 638
rect 1654 542 1657 638
rect 1670 592 1673 718
rect 1806 702 1809 748
rect 1846 712 1849 748
rect 1814 672 1817 708
rect 1694 662 1697 668
rect 1822 662 1825 698
rect 1854 662 1857 848
rect 1902 832 1905 858
rect 1918 852 1921 1058
rect 1946 1048 1950 1051
rect 1930 918 1934 921
rect 1966 882 1969 1058
rect 1998 1052 2001 1068
rect 2022 1052 2025 1158
rect 2046 1052 2049 1068
rect 2022 1032 2025 1048
rect 2026 1018 2030 1021
rect 2006 952 2009 958
rect 1982 942 1985 948
rect 1926 862 1929 868
rect 1946 858 1950 861
rect 1934 852 1937 858
rect 1910 792 1913 838
rect 1954 748 1958 751
rect 1862 742 1865 748
rect 1918 732 1921 738
rect 1926 731 1929 748
rect 1938 738 1942 741
rect 1926 728 1937 731
rect 1870 672 1873 698
rect 1934 692 1937 728
rect 1878 682 1881 688
rect 1914 668 1918 671
rect 1862 662 1865 668
rect 1926 662 1929 668
rect 1682 658 1686 661
rect 1682 648 1686 651
rect 1694 552 1697 558
rect 1734 552 1737 658
rect 1750 642 1753 658
rect 1758 652 1761 658
rect 1766 592 1769 618
rect 1774 562 1777 648
rect 1846 642 1849 658
rect 1614 462 1617 488
rect 1622 402 1625 468
rect 1646 452 1649 458
rect 1622 352 1625 378
rect 1466 178 1470 181
rect 1414 152 1417 168
rect 1422 141 1425 178
rect 1486 172 1489 258
rect 1528 203 1530 207
rect 1534 203 1537 207
rect 1541 203 1544 207
rect 1462 152 1465 168
rect 1550 152 1553 338
rect 1574 292 1577 298
rect 1614 282 1617 308
rect 1630 282 1633 388
rect 1646 292 1649 438
rect 1654 432 1657 538
rect 1662 532 1665 547
rect 1702 542 1705 548
rect 1714 528 1718 531
rect 1742 512 1745 548
rect 1750 532 1753 538
rect 1670 492 1673 508
rect 1670 472 1673 488
rect 1678 472 1681 478
rect 1670 392 1673 458
rect 1678 452 1681 468
rect 1702 452 1705 498
rect 1726 472 1729 488
rect 1774 462 1777 558
rect 1830 551 1833 618
rect 1790 542 1793 548
rect 1798 542 1801 548
rect 1854 541 1857 658
rect 1862 552 1865 658
rect 1890 648 1894 651
rect 1894 622 1897 648
rect 1910 642 1913 658
rect 1918 652 1921 658
rect 1910 592 1913 638
rect 1926 592 1929 628
rect 1922 558 1926 561
rect 1854 538 1865 541
rect 1814 521 1817 538
rect 1806 518 1817 521
rect 1782 462 1785 478
rect 1806 462 1809 518
rect 1846 462 1849 538
rect 1862 462 1865 538
rect 1882 478 1886 481
rect 1902 472 1905 548
rect 1918 502 1921 558
rect 1942 552 1945 738
rect 1954 728 1958 731
rect 1950 682 1953 688
rect 1966 682 1969 878
rect 2014 872 2017 928
rect 2010 858 2014 861
rect 2002 748 2006 751
rect 2022 742 2025 868
rect 1974 702 1977 728
rect 1974 681 1977 698
rect 1990 692 1993 728
rect 1974 678 1982 681
rect 1970 668 1974 671
rect 1962 658 1966 661
rect 1950 622 1953 648
rect 1990 552 1993 678
rect 1998 662 2001 738
rect 2006 682 2009 688
rect 2014 682 2017 688
rect 2022 662 2025 668
rect 2030 662 2033 668
rect 2002 558 2006 561
rect 2038 561 2041 828
rect 2038 558 2049 561
rect 2046 552 2049 558
rect 1930 548 1934 551
rect 1970 548 1974 551
rect 1942 542 1945 548
rect 2038 542 2041 548
rect 1930 538 1934 541
rect 2042 538 2049 541
rect 1902 462 1905 468
rect 1850 458 1854 461
rect 1874 458 1878 461
rect 1682 418 1686 421
rect 1706 418 1710 421
rect 1738 418 1742 421
rect 1734 412 1737 418
rect 1662 332 1665 338
rect 1678 332 1681 398
rect 1694 352 1697 378
rect 1718 342 1721 378
rect 1734 352 1737 368
rect 1786 358 1790 361
rect 1742 352 1745 358
rect 1806 352 1809 458
rect 1862 422 1865 458
rect 1918 432 1921 468
rect 1814 352 1817 368
rect 1678 292 1681 328
rect 1594 278 1598 281
rect 1630 272 1633 278
rect 1670 272 1673 278
rect 1562 268 1566 271
rect 1606 262 1609 268
rect 1642 258 1646 261
rect 1678 261 1681 278
rect 1674 258 1681 261
rect 1558 172 1561 258
rect 1414 138 1425 141
rect 1430 142 1433 148
rect 1414 132 1417 138
rect 1438 72 1441 148
rect 1458 138 1462 141
rect 1446 122 1449 128
rect 1502 72 1505 148
rect 1510 132 1513 148
rect 1566 132 1569 258
rect 1622 252 1625 258
rect 1642 248 1646 251
rect 1598 152 1601 178
rect 1598 142 1601 148
rect 1622 142 1625 178
rect 1630 152 1633 168
rect 1638 132 1641 188
rect 1654 152 1657 158
rect 1654 142 1657 148
rect 1678 142 1681 248
rect 1694 242 1697 338
rect 1726 322 1729 348
rect 1714 318 1721 321
rect 1718 262 1721 318
rect 1686 152 1689 168
rect 1734 152 1737 348
rect 1766 322 1769 348
rect 1774 342 1777 348
rect 1790 332 1793 338
rect 1798 321 1801 328
rect 1790 318 1801 321
rect 1790 292 1793 318
rect 1790 282 1793 288
rect 1806 272 1809 348
rect 1838 342 1841 368
rect 1846 352 1849 418
rect 1894 352 1897 358
rect 1850 348 1857 351
rect 1846 332 1849 338
rect 1814 272 1817 318
rect 1758 262 1761 268
rect 1806 262 1809 268
rect 1758 152 1761 258
rect 1782 152 1785 178
rect 1694 142 1697 148
rect 1566 92 1569 128
rect 1614 92 1617 118
rect 1530 88 1534 91
rect 1590 63 1593 88
rect 1622 82 1625 98
rect 1630 92 1633 128
rect 1638 92 1641 128
rect 1606 72 1609 78
rect 1218 58 1222 61
rect 1670 61 1673 118
rect 1734 92 1737 108
rect 1758 101 1761 148
rect 1806 142 1809 178
rect 1814 152 1817 268
rect 1830 262 1833 318
rect 1822 132 1825 228
rect 1854 172 1857 348
rect 1886 342 1889 348
rect 1870 262 1873 298
rect 1918 292 1921 418
rect 1942 372 1945 538
rect 1950 392 1953 478
rect 1958 462 1961 518
rect 1990 472 1993 528
rect 2006 472 2009 518
rect 2014 512 2017 538
rect 2026 528 2030 531
rect 2034 518 2041 521
rect 2014 492 2017 498
rect 2026 478 2030 481
rect 2026 468 2030 471
rect 2038 462 2041 518
rect 2046 462 2049 538
rect 1930 278 1934 281
rect 1946 278 1953 281
rect 1878 262 1881 278
rect 1902 262 1905 268
rect 1926 262 1929 268
rect 1942 252 1945 258
rect 1894 191 1897 218
rect 1950 192 1953 278
rect 1958 262 1961 388
rect 1982 352 1985 438
rect 1958 222 1961 258
rect 1966 201 1969 218
rect 1958 198 1969 201
rect 1894 188 1905 191
rect 1870 152 1873 168
rect 1834 148 1838 151
rect 1902 151 1905 188
rect 1862 142 1865 148
rect 1826 128 1833 131
rect 1766 112 1769 128
rect 1758 98 1769 101
rect 1718 72 1721 78
rect 1766 72 1769 98
rect 1766 62 1769 68
rect 1798 63 1801 118
rect 1830 92 1833 128
rect 1858 118 1862 121
rect 1670 58 1678 61
rect 1862 62 1865 68
rect 1870 62 1873 118
rect 1886 72 1889 138
rect 1958 62 1961 198
rect 1966 182 1969 188
rect 1974 152 1977 308
rect 1982 262 1985 268
rect 1982 92 1985 258
rect 1990 191 1993 218
rect 1998 202 2001 218
rect 1990 188 1998 191
rect 2006 152 2009 458
rect 2014 351 2017 458
rect 2014 262 2017 328
rect 2026 258 2030 261
rect 1990 102 1993 118
rect 2006 72 2009 128
rect 486 52 489 58
rect 678 52 681 58
rect 1158 52 1161 58
rect 1206 52 1209 58
rect 1270 52 1273 58
rect 658 48 662 51
rect 786 48 790 51
rect 1130 48 1134 51
rect 414 42 417 48
rect 2014 21 2017 98
rect 2026 88 2030 91
rect 2022 62 2025 68
rect 2014 18 2025 21
rect 496 3 498 7
rect 502 3 505 7
rect 509 3 512 7
rect 1528 3 1530 7
rect 1534 3 1537 7
rect 1541 3 1544 7
rect 1990 -18 1993 8
rect 2014 -18 2017 8
rect 1990 -22 1994 -18
rect 2014 -22 2018 -18
rect 2022 -29 2025 18
rect 2030 -19 2034 -18
rect 2038 -19 2041 118
rect 2046 -9 2049 218
rect 2046 -12 2057 -9
rect 2030 -22 2041 -19
rect 2046 -22 2050 -18
rect 2054 -19 2057 -12
rect 2062 -19 2066 -18
rect 2054 -22 2066 -19
rect 2046 -29 2049 -22
rect 2022 -32 2049 -29
<< m3contact >>
rect 498 1803 502 1807
rect 505 1803 509 1807
rect 1530 1803 1534 1807
rect 1537 1803 1541 1807
rect 174 1798 178 1802
rect 814 1798 818 1802
rect 830 1798 834 1802
rect 14 1788 18 1792
rect 54 1788 58 1792
rect 118 1788 122 1792
rect 30 1778 34 1782
rect 6 1578 10 1582
rect 126 1758 130 1762
rect 150 1748 154 1752
rect 606 1748 610 1752
rect 670 1748 674 1752
rect 798 1748 802 1752
rect 94 1688 98 1692
rect 142 1698 146 1702
rect 190 1698 194 1702
rect 166 1688 170 1692
rect 302 1698 306 1702
rect 110 1678 114 1682
rect 286 1678 290 1682
rect 54 1588 58 1592
rect 46 1558 50 1562
rect 30 1548 34 1552
rect 38 1548 42 1552
rect 38 1468 42 1472
rect 166 1658 170 1662
rect 230 1658 234 1662
rect 350 1738 354 1742
rect 374 1738 378 1742
rect 358 1688 362 1692
rect 406 1728 410 1732
rect 446 1718 450 1722
rect 534 1718 538 1722
rect 494 1708 498 1712
rect 510 1708 514 1712
rect 398 1668 402 1672
rect 286 1638 290 1642
rect 174 1548 178 1552
rect 214 1548 218 1552
rect 134 1528 138 1532
rect 166 1528 170 1532
rect 110 1508 114 1512
rect 102 1488 106 1492
rect 94 1478 98 1482
rect 150 1498 154 1502
rect 142 1488 146 1492
rect 166 1478 170 1482
rect 350 1648 354 1652
rect 438 1558 442 1562
rect 278 1488 282 1492
rect 262 1478 266 1482
rect 110 1468 114 1472
rect 126 1468 130 1472
rect 174 1468 178 1472
rect 190 1468 194 1472
rect 246 1468 250 1472
rect 118 1458 122 1462
rect 142 1458 146 1462
rect 182 1458 186 1462
rect 134 1448 138 1452
rect 102 1438 106 1442
rect 94 1338 98 1342
rect 30 1328 34 1332
rect 110 1308 114 1312
rect 110 1288 114 1292
rect 54 1268 58 1272
rect 118 1268 122 1272
rect 134 1258 138 1262
rect 110 1148 114 1152
rect 30 1138 34 1142
rect 54 1088 58 1092
rect 6 1078 10 1082
rect 214 1448 218 1452
rect 206 1438 210 1442
rect 198 1418 202 1422
rect 182 1348 186 1352
rect 206 1388 210 1392
rect 158 1338 162 1342
rect 150 1298 154 1302
rect 302 1418 306 1422
rect 254 1338 258 1342
rect 230 1328 234 1332
rect 294 1318 298 1322
rect 270 1288 274 1292
rect 294 1288 298 1292
rect 150 1278 154 1282
rect 198 1278 202 1282
rect 254 1268 258 1272
rect 158 1248 162 1252
rect 286 1278 290 1282
rect 214 1258 218 1262
rect 246 1258 250 1262
rect 262 1258 266 1262
rect 198 1248 202 1252
rect 142 1128 146 1132
rect 126 1068 130 1072
rect 222 1158 226 1162
rect 278 1248 282 1252
rect 206 1148 210 1152
rect 270 1148 274 1152
rect 166 1098 170 1102
rect 182 1088 186 1092
rect 174 1078 178 1082
rect 230 1128 234 1132
rect 222 1088 226 1092
rect 262 1078 266 1082
rect 278 1078 282 1082
rect 246 1068 250 1072
rect 134 1058 138 1062
rect 150 1058 154 1062
rect 70 1048 74 1052
rect 110 1038 114 1042
rect 126 1038 130 1042
rect 6 988 10 992
rect 126 948 130 952
rect 6 878 10 882
rect 214 1048 218 1052
rect 206 1028 210 1032
rect 182 958 186 962
rect 230 958 234 962
rect 198 948 202 952
rect 206 948 210 952
rect 158 938 162 942
rect 150 898 154 902
rect 206 918 210 922
rect 198 898 202 902
rect 150 888 154 892
rect 174 888 178 892
rect 102 878 106 882
rect 70 868 74 872
rect 86 868 90 872
rect 118 858 122 862
rect 94 818 98 822
rect 118 808 122 812
rect 142 808 146 812
rect 182 878 186 882
rect 190 878 194 882
rect 158 858 162 862
rect 174 858 178 862
rect 158 828 162 832
rect 182 828 186 832
rect 54 748 58 752
rect 134 748 138 752
rect 142 748 146 752
rect 166 748 170 752
rect 118 738 122 742
rect 182 728 186 732
rect 150 708 154 712
rect 102 688 106 692
rect 150 688 154 692
rect 102 668 106 672
rect 142 668 146 672
rect 54 658 58 662
rect 118 658 122 662
rect 62 648 66 652
rect 30 538 34 542
rect 14 468 18 472
rect 14 348 18 352
rect 38 508 42 512
rect 134 658 138 662
rect 150 658 154 662
rect 94 608 98 612
rect 126 588 130 592
rect 110 528 114 532
rect 78 518 82 522
rect 86 518 90 522
rect 110 508 114 512
rect 142 568 146 572
rect 134 538 138 542
rect 94 468 98 472
rect 126 468 130 472
rect 118 458 122 462
rect 118 388 122 392
rect 54 368 58 372
rect 190 678 194 682
rect 182 658 186 662
rect 166 648 170 652
rect 182 558 186 562
rect 150 458 154 462
rect 134 388 138 392
rect 214 908 218 912
rect 310 1278 314 1282
rect 310 1268 314 1272
rect 518 1658 522 1662
rect 534 1658 538 1662
rect 462 1628 466 1632
rect 498 1603 502 1607
rect 505 1603 509 1607
rect 574 1708 578 1712
rect 918 1788 922 1792
rect 1950 1758 1954 1762
rect 918 1748 922 1752
rect 1214 1748 1218 1752
rect 1934 1748 1938 1752
rect 654 1738 658 1742
rect 774 1738 778 1742
rect 854 1738 858 1742
rect 910 1738 914 1742
rect 942 1738 946 1742
rect 1006 1738 1010 1742
rect 662 1728 666 1732
rect 574 1668 578 1672
rect 582 1648 586 1652
rect 590 1618 594 1622
rect 614 1618 618 1622
rect 550 1598 554 1602
rect 526 1568 530 1572
rect 526 1548 530 1552
rect 358 1528 362 1532
rect 382 1528 386 1532
rect 358 1478 362 1482
rect 494 1478 498 1482
rect 446 1468 450 1472
rect 462 1468 466 1472
rect 382 1358 386 1362
rect 390 1288 394 1292
rect 350 1258 354 1262
rect 366 1258 370 1262
rect 374 1248 378 1252
rect 646 1658 650 1662
rect 630 1588 634 1592
rect 574 1558 578 1562
rect 614 1558 618 1562
rect 630 1558 634 1562
rect 566 1548 570 1552
rect 598 1548 602 1552
rect 558 1498 562 1502
rect 542 1478 546 1482
rect 550 1478 554 1482
rect 590 1538 594 1542
rect 598 1518 602 1522
rect 630 1488 634 1492
rect 686 1718 690 1722
rect 678 1658 682 1662
rect 646 1538 650 1542
rect 558 1468 562 1472
rect 574 1468 578 1472
rect 582 1468 586 1472
rect 638 1468 642 1472
rect 518 1458 522 1462
rect 518 1448 522 1452
rect 542 1448 546 1452
rect 654 1518 658 1522
rect 670 1508 674 1512
rect 662 1478 666 1482
rect 598 1448 602 1452
rect 590 1438 594 1442
rect 558 1428 562 1432
rect 582 1428 586 1432
rect 498 1403 502 1407
rect 505 1403 509 1407
rect 462 1368 466 1372
rect 422 1348 426 1352
rect 414 1338 418 1342
rect 406 1328 410 1332
rect 422 1328 426 1332
rect 430 1308 434 1312
rect 470 1348 474 1352
rect 494 1348 498 1352
rect 526 1368 530 1372
rect 566 1348 570 1352
rect 478 1338 482 1342
rect 454 1328 458 1332
rect 446 1318 450 1322
rect 446 1308 450 1312
rect 446 1298 450 1302
rect 430 1288 434 1292
rect 438 1288 442 1292
rect 406 1258 410 1262
rect 438 1278 442 1282
rect 398 1178 402 1182
rect 302 1148 306 1152
rect 454 1288 458 1292
rect 558 1328 562 1332
rect 526 1318 530 1322
rect 470 1278 474 1282
rect 494 1298 498 1302
rect 502 1278 506 1282
rect 478 1268 482 1272
rect 486 1268 490 1272
rect 510 1258 514 1262
rect 462 1238 466 1242
rect 446 1228 450 1232
rect 478 1228 482 1232
rect 494 1228 498 1232
rect 438 1218 442 1222
rect 430 1168 434 1172
rect 422 1158 426 1162
rect 382 1148 386 1152
rect 414 1148 418 1152
rect 438 1148 442 1152
rect 374 1128 378 1132
rect 422 1138 426 1142
rect 406 1128 410 1132
rect 398 1098 402 1102
rect 470 1218 474 1222
rect 462 1178 466 1182
rect 498 1203 502 1207
rect 505 1203 509 1207
rect 638 1338 642 1342
rect 598 1318 602 1322
rect 558 1308 562 1312
rect 574 1288 578 1292
rect 598 1278 602 1282
rect 606 1278 610 1282
rect 590 1268 594 1272
rect 654 1358 658 1362
rect 662 1358 666 1362
rect 678 1408 682 1412
rect 710 1718 714 1722
rect 822 1718 826 1722
rect 822 1708 826 1712
rect 814 1668 818 1672
rect 902 1668 906 1672
rect 710 1618 714 1622
rect 710 1558 714 1562
rect 790 1648 794 1652
rect 926 1728 930 1732
rect 1018 1703 1022 1707
rect 1025 1703 1029 1707
rect 974 1688 978 1692
rect 990 1688 994 1692
rect 1142 1738 1146 1742
rect 1350 1738 1354 1742
rect 1390 1738 1394 1742
rect 1462 1738 1466 1742
rect 1486 1738 1490 1742
rect 1510 1738 1514 1742
rect 1574 1738 1578 1742
rect 1150 1728 1154 1732
rect 1214 1728 1218 1732
rect 1230 1728 1234 1732
rect 1294 1728 1298 1732
rect 1118 1718 1122 1722
rect 1190 1718 1194 1722
rect 990 1678 994 1682
rect 1006 1678 1010 1682
rect 1094 1678 1098 1682
rect 1046 1668 1050 1672
rect 1070 1668 1074 1672
rect 1158 1668 1162 1672
rect 1174 1668 1178 1672
rect 942 1648 946 1652
rect 758 1618 762 1622
rect 798 1618 802 1622
rect 822 1618 826 1622
rect 750 1608 754 1612
rect 742 1558 746 1562
rect 782 1608 786 1612
rect 838 1588 842 1592
rect 758 1568 762 1572
rect 774 1568 778 1572
rect 846 1548 850 1552
rect 774 1538 778 1542
rect 694 1508 698 1512
rect 750 1508 754 1512
rect 718 1498 722 1502
rect 758 1488 762 1492
rect 702 1378 706 1382
rect 686 1358 690 1362
rect 734 1358 738 1362
rect 702 1348 706 1352
rect 982 1638 986 1642
rect 974 1578 978 1582
rect 1030 1608 1034 1612
rect 958 1538 962 1542
rect 1006 1538 1010 1542
rect 1046 1538 1050 1542
rect 862 1488 866 1492
rect 950 1488 954 1492
rect 838 1478 842 1482
rect 862 1468 866 1472
rect 894 1468 898 1472
rect 782 1398 786 1402
rect 806 1398 810 1402
rect 742 1348 746 1352
rect 774 1348 778 1352
rect 790 1348 794 1352
rect 662 1338 666 1342
rect 694 1338 698 1342
rect 710 1338 714 1342
rect 678 1318 682 1322
rect 678 1278 682 1282
rect 702 1288 706 1292
rect 670 1268 674 1272
rect 702 1268 706 1272
rect 542 1248 546 1252
rect 534 1238 538 1242
rect 558 1238 562 1242
rect 630 1228 634 1232
rect 550 1218 554 1222
rect 614 1188 618 1192
rect 582 1178 586 1182
rect 534 1158 538 1162
rect 470 1138 474 1142
rect 486 1138 490 1142
rect 454 1108 458 1112
rect 478 1128 482 1132
rect 470 1098 474 1102
rect 358 1088 362 1092
rect 318 1078 322 1082
rect 302 1068 306 1072
rect 350 1068 354 1072
rect 270 1058 274 1062
rect 326 1058 330 1062
rect 406 1078 410 1082
rect 438 1078 442 1082
rect 462 1078 466 1082
rect 470 1078 474 1082
rect 662 1258 666 1262
rect 678 1248 682 1252
rect 710 1248 714 1252
rect 654 1238 658 1242
rect 638 1188 642 1192
rect 638 1178 642 1182
rect 518 1138 522 1142
rect 558 1138 562 1142
rect 606 1138 610 1142
rect 638 1138 642 1142
rect 526 1128 530 1132
rect 614 1128 618 1132
rect 638 1128 642 1132
rect 550 1108 554 1112
rect 550 1098 554 1102
rect 582 1098 586 1102
rect 574 1088 578 1092
rect 374 1068 378 1072
rect 422 1068 426 1072
rect 454 1068 458 1072
rect 510 1068 514 1072
rect 518 1058 522 1062
rect 526 1058 530 1062
rect 574 1058 578 1062
rect 270 1038 274 1042
rect 334 1038 338 1042
rect 374 1028 378 1032
rect 278 988 282 992
rect 302 968 306 972
rect 318 948 322 952
rect 334 948 338 952
rect 366 968 370 972
rect 422 1048 426 1052
rect 430 1048 434 1052
rect 398 1038 402 1042
rect 382 988 386 992
rect 498 1003 502 1007
rect 505 1003 509 1007
rect 478 988 482 992
rect 478 978 482 982
rect 414 958 418 962
rect 454 958 458 962
rect 270 928 274 932
rect 286 928 290 932
rect 278 908 282 912
rect 254 888 258 892
rect 230 878 234 882
rect 254 878 258 882
rect 278 878 282 882
rect 222 858 226 862
rect 238 798 242 802
rect 222 788 226 792
rect 270 788 274 792
rect 214 758 218 762
rect 294 908 298 912
rect 334 938 338 942
rect 358 928 362 932
rect 398 928 402 932
rect 302 898 306 902
rect 310 898 314 902
rect 342 898 346 902
rect 374 898 378 902
rect 374 888 378 892
rect 358 868 362 872
rect 390 868 394 872
rect 342 858 346 862
rect 310 798 314 802
rect 302 768 306 772
rect 246 738 250 742
rect 246 698 250 702
rect 286 698 290 702
rect 270 678 274 682
rect 278 678 282 682
rect 294 678 298 682
rect 262 668 266 672
rect 254 658 258 662
rect 334 748 338 752
rect 366 748 370 752
rect 350 728 354 732
rect 318 718 322 722
rect 334 678 338 682
rect 302 668 306 672
rect 302 658 306 662
rect 326 658 330 662
rect 286 648 290 652
rect 246 578 250 582
rect 214 568 218 572
rect 198 558 202 562
rect 222 558 226 562
rect 190 548 194 552
rect 246 548 250 552
rect 198 538 202 542
rect 166 458 170 462
rect 182 448 186 452
rect 190 438 194 442
rect 238 488 242 492
rect 222 458 226 462
rect 230 448 234 452
rect 222 438 226 442
rect 158 368 162 372
rect 198 368 202 372
rect 158 358 162 362
rect 182 358 186 362
rect 142 348 146 352
rect 102 328 106 332
rect 70 318 74 322
rect 62 258 66 262
rect 174 338 178 342
rect 190 338 194 342
rect 158 328 162 332
rect 126 318 130 322
rect 166 318 170 322
rect 198 318 202 322
rect 134 268 138 272
rect 150 228 154 232
rect 102 158 106 162
rect 118 158 122 162
rect 110 148 114 152
rect 142 148 146 152
rect 54 128 58 132
rect 278 459 282 463
rect 326 648 330 652
rect 310 638 314 642
rect 326 638 330 642
rect 302 618 306 622
rect 374 658 378 662
rect 406 858 410 862
rect 398 848 402 852
rect 390 838 394 842
rect 422 928 426 932
rect 422 918 426 922
rect 430 898 434 902
rect 494 968 498 972
rect 454 938 458 942
rect 486 938 490 942
rect 446 918 450 922
rect 438 888 442 892
rect 454 888 458 892
rect 502 888 506 892
rect 438 878 442 882
rect 414 818 418 822
rect 454 858 458 862
rect 422 798 426 802
rect 566 1038 570 1042
rect 558 1028 562 1032
rect 582 1018 586 1022
rect 606 1008 610 1012
rect 582 968 586 972
rect 550 948 554 952
rect 534 938 538 942
rect 574 938 578 942
rect 590 938 594 942
rect 678 1228 682 1232
rect 758 1318 762 1322
rect 806 1318 810 1322
rect 814 1318 818 1322
rect 766 1308 770 1312
rect 782 1308 786 1312
rect 766 1258 770 1262
rect 758 1248 762 1252
rect 742 1238 746 1242
rect 822 1298 826 1302
rect 838 1278 842 1282
rect 854 1278 858 1282
rect 958 1468 962 1472
rect 1018 1503 1022 1507
rect 1025 1503 1029 1507
rect 1046 1468 1050 1472
rect 998 1458 1002 1462
rect 870 1428 874 1432
rect 894 1428 898 1432
rect 1222 1718 1226 1722
rect 1262 1698 1266 1702
rect 1246 1678 1250 1682
rect 1254 1678 1258 1682
rect 1246 1668 1250 1672
rect 1254 1668 1258 1672
rect 1110 1658 1114 1662
rect 1142 1658 1146 1662
rect 1182 1658 1186 1662
rect 1206 1658 1210 1662
rect 1062 1638 1066 1642
rect 1086 1638 1090 1642
rect 1070 1628 1074 1632
rect 1086 1568 1090 1572
rect 1070 1548 1074 1552
rect 1118 1648 1122 1652
rect 1126 1578 1130 1582
rect 1214 1648 1218 1652
rect 1254 1648 1258 1652
rect 1174 1638 1178 1642
rect 1206 1638 1210 1642
rect 1166 1628 1170 1632
rect 1150 1618 1154 1622
rect 1142 1568 1146 1572
rect 1150 1568 1154 1572
rect 1126 1548 1130 1552
rect 1102 1538 1106 1542
rect 1134 1538 1138 1542
rect 1094 1518 1098 1522
rect 1110 1518 1114 1522
rect 1070 1508 1074 1512
rect 1118 1498 1122 1502
rect 1118 1468 1122 1472
rect 1166 1578 1170 1582
rect 1174 1568 1178 1572
rect 1158 1558 1162 1562
rect 1150 1538 1154 1542
rect 1038 1458 1042 1462
rect 1062 1458 1066 1462
rect 1190 1558 1194 1562
rect 1190 1518 1194 1522
rect 1198 1508 1202 1512
rect 1230 1608 1234 1612
rect 1214 1588 1218 1592
rect 1246 1588 1250 1592
rect 1214 1538 1218 1542
rect 1230 1518 1234 1522
rect 1238 1508 1242 1512
rect 1190 1478 1194 1482
rect 1206 1478 1210 1482
rect 1214 1478 1218 1482
rect 1182 1468 1186 1472
rect 1022 1448 1026 1452
rect 1150 1448 1154 1452
rect 1174 1448 1178 1452
rect 1102 1438 1106 1442
rect 1174 1438 1178 1442
rect 1070 1428 1074 1432
rect 1038 1398 1042 1402
rect 1078 1398 1082 1402
rect 1094 1388 1098 1392
rect 1038 1378 1042 1382
rect 1054 1378 1058 1382
rect 918 1368 922 1372
rect 1014 1368 1018 1372
rect 886 1358 890 1362
rect 1022 1358 1026 1362
rect 942 1348 946 1352
rect 934 1338 938 1342
rect 870 1308 874 1312
rect 926 1308 930 1312
rect 870 1298 874 1302
rect 918 1298 922 1302
rect 902 1288 906 1292
rect 886 1278 890 1282
rect 862 1268 866 1272
rect 806 1258 810 1262
rect 830 1248 834 1252
rect 862 1258 866 1262
rect 942 1258 946 1262
rect 846 1238 850 1242
rect 862 1238 866 1242
rect 782 1228 786 1232
rect 790 1228 794 1232
rect 750 1218 754 1222
rect 686 1208 690 1212
rect 654 1118 658 1122
rect 678 1118 682 1122
rect 646 1098 650 1102
rect 670 1098 674 1102
rect 646 1088 650 1092
rect 702 1108 706 1112
rect 718 1098 722 1102
rect 702 1088 706 1092
rect 694 1078 698 1082
rect 670 1068 674 1072
rect 622 998 626 1002
rect 646 998 650 1002
rect 718 1078 722 1082
rect 766 1148 770 1152
rect 694 1058 698 1062
rect 726 1058 730 1062
rect 678 1048 682 1052
rect 654 968 658 972
rect 662 948 666 952
rect 646 938 650 942
rect 598 918 602 922
rect 646 918 650 922
rect 558 908 562 912
rect 614 908 618 912
rect 590 888 594 892
rect 638 888 642 892
rect 630 878 634 882
rect 550 859 554 863
rect 670 908 674 912
rect 662 898 666 902
rect 694 1038 698 1042
rect 766 1128 770 1132
rect 838 1188 842 1192
rect 798 1148 802 1152
rect 822 1118 826 1122
rect 750 1068 754 1072
rect 734 1018 738 1022
rect 718 998 722 1002
rect 718 988 722 992
rect 758 1008 762 1012
rect 742 978 746 982
rect 782 988 786 992
rect 766 968 770 972
rect 822 1098 826 1102
rect 854 1178 858 1182
rect 870 1178 874 1182
rect 862 1158 866 1162
rect 918 1168 922 1172
rect 878 1158 882 1162
rect 862 1148 866 1152
rect 974 1338 978 1342
rect 982 1318 986 1322
rect 1018 1303 1022 1307
rect 1025 1303 1029 1307
rect 990 1288 994 1292
rect 998 1258 1002 1262
rect 1006 1258 1010 1262
rect 966 1158 970 1162
rect 958 1148 962 1152
rect 894 1138 898 1142
rect 830 1088 834 1092
rect 798 1078 802 1082
rect 806 1008 810 1012
rect 790 968 794 972
rect 790 948 794 952
rect 742 938 746 942
rect 686 918 690 922
rect 734 918 738 922
rect 726 908 730 912
rect 718 888 722 892
rect 782 938 786 942
rect 758 928 762 932
rect 742 888 746 892
rect 814 988 818 992
rect 830 968 834 972
rect 830 948 834 952
rect 854 1088 858 1092
rect 878 1088 882 1092
rect 974 1128 978 1132
rect 902 1088 906 1092
rect 942 1088 946 1092
rect 886 1078 890 1082
rect 902 1078 906 1082
rect 894 1068 898 1072
rect 934 1068 938 1072
rect 998 1068 1002 1072
rect 854 1058 858 1062
rect 870 1058 874 1062
rect 966 1058 970 1062
rect 910 1048 914 1052
rect 854 1038 858 1042
rect 902 1038 906 1042
rect 862 968 866 972
rect 854 948 858 952
rect 974 1048 978 1052
rect 918 1038 922 1042
rect 910 1028 914 1032
rect 934 988 938 992
rect 918 978 922 982
rect 750 868 754 872
rect 798 868 802 872
rect 606 858 610 862
rect 614 848 618 852
rect 630 848 634 852
rect 646 828 650 832
rect 654 828 658 832
rect 526 818 530 822
rect 582 818 586 822
rect 498 803 502 807
rect 505 803 509 807
rect 478 798 482 802
rect 454 788 458 792
rect 422 778 426 782
rect 398 768 402 772
rect 382 588 386 592
rect 342 568 346 572
rect 302 548 306 552
rect 326 488 330 492
rect 446 758 450 762
rect 502 788 506 792
rect 486 758 490 762
rect 510 758 514 762
rect 438 748 442 752
rect 470 748 474 752
rect 478 748 482 752
rect 510 748 514 752
rect 462 738 466 742
rect 438 728 442 732
rect 478 728 482 732
rect 462 698 466 702
rect 534 788 538 792
rect 526 778 530 782
rect 550 768 554 772
rect 542 758 546 762
rect 534 738 538 742
rect 518 708 522 712
rect 486 688 490 692
rect 478 678 482 682
rect 502 678 506 682
rect 422 668 426 672
rect 470 668 474 672
rect 510 668 514 672
rect 526 668 530 672
rect 462 658 466 662
rect 422 638 426 642
rect 414 628 418 632
rect 462 638 466 642
rect 446 608 450 612
rect 430 588 434 592
rect 414 578 418 582
rect 374 558 378 562
rect 398 558 402 562
rect 374 548 378 552
rect 390 538 394 542
rect 390 508 394 512
rect 350 478 354 482
rect 390 478 394 482
rect 318 378 322 382
rect 286 358 290 362
rect 326 358 330 362
rect 374 468 378 472
rect 350 458 354 462
rect 374 458 378 462
rect 422 468 426 472
rect 406 418 410 422
rect 382 388 386 392
rect 358 368 362 372
rect 374 368 378 372
rect 278 348 282 352
rect 350 348 354 352
rect 302 338 306 342
rect 230 278 234 282
rect 286 308 290 312
rect 254 268 258 272
rect 222 258 226 262
rect 526 648 530 652
rect 498 603 502 607
rect 505 603 509 607
rect 470 578 474 582
rect 470 568 474 572
rect 510 558 514 562
rect 526 548 530 552
rect 614 778 618 782
rect 606 748 610 752
rect 678 758 682 762
rect 742 858 746 862
rect 774 858 778 862
rect 718 848 722 852
rect 806 848 810 852
rect 726 838 730 842
rect 782 838 786 842
rect 702 808 706 812
rect 726 808 730 812
rect 838 928 842 932
rect 846 928 850 932
rect 822 898 826 902
rect 830 888 834 892
rect 830 868 834 872
rect 838 858 842 862
rect 830 828 834 832
rect 766 788 770 792
rect 806 788 810 792
rect 702 758 706 762
rect 718 758 722 762
rect 630 748 634 752
rect 662 748 666 752
rect 670 748 674 752
rect 838 768 842 772
rect 734 748 738 752
rect 750 748 754 752
rect 758 748 762 752
rect 790 748 794 752
rect 590 738 594 742
rect 622 738 626 742
rect 662 738 666 742
rect 678 738 682 742
rect 710 738 714 742
rect 606 718 610 722
rect 582 698 586 702
rect 590 688 594 692
rect 686 728 690 732
rect 654 688 658 692
rect 710 688 714 692
rect 590 678 594 682
rect 646 678 650 682
rect 550 668 554 672
rect 542 658 546 662
rect 558 648 562 652
rect 566 648 570 652
rect 582 638 586 642
rect 574 578 578 582
rect 566 568 570 572
rect 558 558 562 562
rect 518 488 522 492
rect 534 488 538 492
rect 454 468 458 472
rect 446 458 450 462
rect 438 428 442 432
rect 526 448 530 452
rect 510 418 514 422
rect 498 403 502 407
rect 505 403 509 407
rect 518 378 522 382
rect 398 358 402 362
rect 406 348 410 352
rect 430 358 434 362
rect 462 358 466 362
rect 478 358 482 362
rect 438 338 442 342
rect 486 338 490 342
rect 390 328 394 332
rect 462 328 466 332
rect 334 318 338 322
rect 470 318 474 322
rect 414 298 418 302
rect 510 298 514 302
rect 310 288 314 292
rect 342 288 346 292
rect 462 288 466 292
rect 326 278 330 282
rect 358 278 362 282
rect 438 278 442 282
rect 398 268 402 272
rect 454 268 458 272
rect 326 258 330 262
rect 254 168 258 172
rect 302 168 306 172
rect 318 168 322 172
rect 262 158 266 162
rect 294 158 298 162
rect 198 148 202 152
rect 278 148 282 152
rect 318 148 322 152
rect 382 248 386 252
rect 382 188 386 192
rect 342 168 346 172
rect 494 278 498 282
rect 478 268 482 272
rect 462 258 466 262
rect 486 248 490 252
rect 502 248 506 252
rect 454 238 458 242
rect 498 203 502 207
rect 505 203 509 207
rect 502 178 506 182
rect 518 168 522 172
rect 342 148 346 152
rect 94 138 98 142
rect 150 138 154 142
rect 262 138 266 142
rect 318 138 322 142
rect 326 138 330 142
rect 366 138 370 142
rect 382 138 386 142
rect 446 148 450 152
rect 534 438 538 442
rect 566 528 570 532
rect 582 568 586 572
rect 598 608 602 612
rect 606 588 610 592
rect 598 548 602 552
rect 574 508 578 512
rect 550 448 554 452
rect 566 428 570 432
rect 574 398 578 402
rect 590 508 594 512
rect 606 488 610 492
rect 702 678 706 682
rect 726 678 730 682
rect 702 668 706 672
rect 710 658 714 662
rect 734 648 738 652
rect 782 738 786 742
rect 822 738 826 742
rect 838 738 842 742
rect 758 728 762 732
rect 798 728 802 732
rect 806 728 810 732
rect 830 728 834 732
rect 790 698 794 702
rect 758 688 762 692
rect 750 668 754 672
rect 742 628 746 632
rect 662 618 666 622
rect 622 608 626 612
rect 630 578 634 582
rect 630 568 634 572
rect 622 538 626 542
rect 638 538 642 542
rect 654 538 658 542
rect 710 548 714 552
rect 774 628 778 632
rect 790 598 794 602
rect 766 578 770 582
rect 766 548 770 552
rect 774 548 778 552
rect 798 548 802 552
rect 750 538 754 542
rect 646 478 650 482
rect 766 528 770 532
rect 750 478 754 482
rect 814 658 818 662
rect 814 578 818 582
rect 854 908 858 912
rect 934 948 938 952
rect 894 928 898 932
rect 910 928 914 932
rect 886 908 890 912
rect 870 898 874 902
rect 854 888 858 892
rect 902 888 906 892
rect 878 868 882 872
rect 926 868 930 872
rect 862 838 866 842
rect 862 778 866 782
rect 854 718 858 722
rect 846 668 850 672
rect 982 1038 986 1042
rect 966 948 970 952
rect 910 838 914 842
rect 966 838 970 842
rect 918 818 922 822
rect 942 818 946 822
rect 942 808 946 812
rect 918 768 922 772
rect 934 768 938 772
rect 878 758 882 762
rect 886 758 890 762
rect 894 738 898 742
rect 910 738 914 742
rect 886 718 890 722
rect 902 718 906 722
rect 878 708 882 712
rect 870 688 874 692
rect 870 678 874 682
rect 934 748 938 752
rect 990 978 994 982
rect 990 938 994 942
rect 990 858 994 862
rect 974 798 978 802
rect 1022 1128 1026 1132
rect 1018 1103 1022 1107
rect 1025 1103 1029 1107
rect 1094 1348 1098 1352
rect 1046 1308 1050 1312
rect 1046 1268 1050 1272
rect 1054 1258 1058 1262
rect 1222 1458 1226 1462
rect 1246 1498 1250 1502
rect 1254 1488 1258 1492
rect 1206 1438 1210 1442
rect 1230 1438 1234 1442
rect 1438 1728 1442 1732
rect 1406 1698 1410 1702
rect 1342 1678 1346 1682
rect 1286 1668 1290 1672
rect 1286 1658 1290 1662
rect 1278 1578 1282 1582
rect 1510 1728 1514 1732
rect 1326 1638 1330 1642
rect 1454 1638 1458 1642
rect 1294 1558 1298 1562
rect 1286 1508 1290 1512
rect 1334 1538 1338 1542
rect 1334 1508 1338 1512
rect 1662 1738 1666 1742
rect 1734 1728 1738 1732
rect 1614 1688 1618 1692
rect 1542 1658 1546 1662
rect 1590 1658 1594 1662
rect 1530 1603 1534 1607
rect 1537 1603 1541 1607
rect 1582 1548 1586 1552
rect 1510 1538 1514 1542
rect 1382 1528 1386 1532
rect 1470 1528 1474 1532
rect 1438 1518 1442 1522
rect 1462 1518 1466 1522
rect 1358 1508 1362 1512
rect 1350 1498 1354 1502
rect 1406 1498 1410 1502
rect 1430 1488 1434 1492
rect 1310 1478 1314 1482
rect 1374 1468 1378 1472
rect 1294 1458 1298 1462
rect 1318 1458 1322 1462
rect 1366 1458 1370 1462
rect 1254 1448 1258 1452
rect 1270 1448 1274 1452
rect 1278 1448 1282 1452
rect 1294 1448 1298 1452
rect 1262 1438 1266 1442
rect 1286 1438 1290 1442
rect 1182 1428 1186 1432
rect 1246 1428 1250 1432
rect 1270 1428 1274 1432
rect 1158 1398 1162 1402
rect 1110 1378 1114 1382
rect 1134 1378 1138 1382
rect 1142 1348 1146 1352
rect 1078 1318 1082 1322
rect 1102 1318 1106 1322
rect 1086 1278 1090 1282
rect 1094 1278 1098 1282
rect 1078 1268 1082 1272
rect 1102 1268 1106 1272
rect 1110 1258 1114 1262
rect 1126 1258 1130 1262
rect 1078 1248 1082 1252
rect 1062 1228 1066 1232
rect 1102 1228 1106 1232
rect 1134 1238 1138 1242
rect 1118 1218 1122 1222
rect 1158 1308 1162 1312
rect 1150 1298 1154 1302
rect 1158 1288 1162 1292
rect 1182 1408 1186 1412
rect 1230 1408 1234 1412
rect 1190 1368 1194 1372
rect 1254 1368 1258 1372
rect 1262 1368 1266 1372
rect 1214 1347 1218 1351
rect 1286 1388 1290 1392
rect 1278 1378 1282 1382
rect 1310 1408 1314 1412
rect 1350 1438 1354 1442
rect 1614 1658 1618 1662
rect 1670 1688 1674 1692
rect 1646 1638 1650 1642
rect 1654 1638 1658 1642
rect 1718 1598 1722 1602
rect 1822 1738 1826 1742
rect 1934 1728 1938 1732
rect 1902 1708 1906 1712
rect 1806 1688 1810 1692
rect 1846 1688 1850 1692
rect 1902 1688 1906 1692
rect 1878 1678 1882 1682
rect 1950 1738 1954 1742
rect 2006 1768 2010 1772
rect 2046 1748 2050 1752
rect 2014 1728 2018 1732
rect 2022 1728 2026 1732
rect 1966 1718 1970 1722
rect 1958 1708 1962 1712
rect 2006 1708 2010 1712
rect 1982 1678 1986 1682
rect 1838 1668 1842 1672
rect 1910 1668 1914 1672
rect 1894 1658 1898 1662
rect 1798 1648 1802 1652
rect 1838 1648 1842 1652
rect 1870 1648 1874 1652
rect 1734 1578 1738 1582
rect 1622 1548 1626 1552
rect 1694 1538 1698 1542
rect 1790 1558 1794 1562
rect 1806 1548 1810 1552
rect 1734 1528 1738 1532
rect 1678 1518 1682 1522
rect 1598 1498 1602 1502
rect 1630 1498 1634 1502
rect 1526 1488 1530 1492
rect 1542 1488 1546 1492
rect 1462 1478 1466 1482
rect 1518 1478 1522 1482
rect 1614 1478 1618 1482
rect 1438 1458 1442 1462
rect 1422 1438 1426 1442
rect 1382 1418 1386 1422
rect 1414 1398 1418 1402
rect 1406 1378 1410 1382
rect 1318 1358 1322 1362
rect 1342 1358 1346 1362
rect 1310 1348 1314 1352
rect 1358 1348 1362 1352
rect 1382 1348 1386 1352
rect 1174 1308 1178 1312
rect 1182 1298 1186 1302
rect 1254 1328 1258 1332
rect 1318 1328 1322 1332
rect 1342 1328 1346 1332
rect 1350 1308 1354 1312
rect 1310 1278 1314 1282
rect 1230 1258 1234 1262
rect 1310 1248 1314 1252
rect 1350 1248 1354 1252
rect 1166 1238 1170 1242
rect 1222 1238 1226 1242
rect 1174 1228 1178 1232
rect 1078 1188 1082 1192
rect 1086 1188 1090 1192
rect 1062 1158 1066 1162
rect 1190 1168 1194 1172
rect 1094 1158 1098 1162
rect 1054 1138 1058 1142
rect 1078 1138 1082 1142
rect 1110 1138 1114 1142
rect 1182 1138 1186 1142
rect 1046 1068 1050 1072
rect 1022 1058 1026 1062
rect 1030 1048 1034 1052
rect 1022 1008 1026 1012
rect 1018 903 1022 907
rect 1025 903 1029 907
rect 1046 1038 1050 1042
rect 1078 968 1082 972
rect 1126 1118 1130 1122
rect 1150 1118 1154 1122
rect 1134 1078 1138 1082
rect 1206 1158 1210 1162
rect 1206 1118 1210 1122
rect 1214 1088 1218 1092
rect 1206 1068 1210 1072
rect 1102 1058 1106 1062
rect 1142 1028 1146 1032
rect 1054 948 1058 952
rect 1086 948 1090 952
rect 1134 948 1138 952
rect 1054 888 1058 892
rect 1006 878 1010 882
rect 1038 878 1042 882
rect 1174 1028 1178 1032
rect 1150 978 1154 982
rect 1166 978 1170 982
rect 1182 968 1186 972
rect 1158 948 1162 952
rect 1126 938 1130 942
rect 1006 858 1010 862
rect 1038 858 1042 862
rect 1062 858 1066 862
rect 1030 848 1034 852
rect 998 778 1002 782
rect 958 768 962 772
rect 1102 848 1106 852
rect 974 758 978 762
rect 1046 758 1050 762
rect 1086 758 1090 762
rect 1118 758 1122 762
rect 966 748 970 752
rect 974 738 978 742
rect 950 728 954 732
rect 990 688 994 692
rect 934 668 938 672
rect 990 668 994 672
rect 902 658 906 662
rect 934 658 938 662
rect 838 648 842 652
rect 830 568 834 572
rect 966 648 970 652
rect 846 638 850 642
rect 862 638 866 642
rect 854 628 858 632
rect 846 568 850 572
rect 878 618 882 622
rect 886 608 890 612
rect 870 598 874 602
rect 774 468 778 472
rect 614 458 618 462
rect 710 458 714 462
rect 614 378 618 382
rect 558 358 562 362
rect 598 358 602 362
rect 750 438 754 442
rect 694 428 698 432
rect 686 388 690 392
rect 638 358 642 362
rect 646 358 650 362
rect 654 358 658 362
rect 670 358 674 362
rect 654 348 658 352
rect 534 338 538 342
rect 582 338 586 342
rect 662 338 666 342
rect 686 338 690 342
rect 750 408 754 412
rect 734 398 738 402
rect 806 468 810 472
rect 806 368 810 372
rect 750 358 754 362
rect 574 328 578 332
rect 542 308 546 312
rect 550 298 554 302
rect 558 268 562 272
rect 550 258 554 262
rect 590 308 594 312
rect 614 298 618 302
rect 590 258 594 262
rect 614 268 618 272
rect 694 318 698 322
rect 670 298 674 302
rect 630 278 634 282
rect 718 298 722 302
rect 830 518 834 522
rect 838 518 842 522
rect 982 598 986 602
rect 894 558 898 562
rect 910 558 914 562
rect 926 558 930 562
rect 966 558 970 562
rect 870 528 874 532
rect 878 528 882 532
rect 902 528 906 532
rect 934 528 938 532
rect 838 508 842 512
rect 846 508 850 512
rect 886 508 890 512
rect 822 478 826 482
rect 830 478 834 482
rect 822 448 826 452
rect 822 408 826 412
rect 830 398 834 402
rect 774 348 778 352
rect 758 328 762 332
rect 798 328 802 332
rect 654 268 658 272
rect 694 268 698 272
rect 718 268 722 272
rect 630 248 634 252
rect 654 238 658 242
rect 598 228 602 232
rect 606 228 610 232
rect 622 228 626 232
rect 566 178 570 182
rect 550 168 554 172
rect 622 218 626 222
rect 662 218 666 222
rect 734 258 738 262
rect 726 248 730 252
rect 742 248 746 252
rect 686 228 690 232
rect 678 188 682 192
rect 678 168 682 172
rect 614 148 618 152
rect 430 138 434 142
rect 534 138 538 142
rect 110 128 114 132
rect 358 128 362 132
rect 390 128 394 132
rect 398 128 402 132
rect 414 128 418 132
rect 390 118 394 122
rect 262 108 266 112
rect 286 108 290 112
rect 246 98 250 102
rect 14 68 18 72
rect 70 68 74 72
rect 142 58 146 62
rect 158 58 162 62
rect 190 58 194 62
rect 270 58 274 62
rect 286 58 290 62
rect 310 58 314 62
rect 414 88 418 92
rect 574 118 578 122
rect 598 68 602 72
rect 702 238 706 242
rect 694 188 698 192
rect 726 168 730 172
rect 870 498 874 502
rect 878 488 882 492
rect 846 468 850 472
rect 918 508 922 512
rect 910 488 914 492
rect 958 498 962 502
rect 950 488 954 492
rect 926 468 930 472
rect 950 468 954 472
rect 846 388 850 392
rect 862 448 866 452
rect 1158 928 1162 932
rect 1158 888 1162 892
rect 1174 948 1178 952
rect 1230 1218 1234 1222
rect 1238 1198 1242 1202
rect 1294 1168 1298 1172
rect 1302 1148 1306 1152
rect 1326 1168 1330 1172
rect 1254 1138 1258 1142
rect 1294 1138 1298 1142
rect 1318 1138 1322 1142
rect 1246 1108 1250 1112
rect 1238 1098 1242 1102
rect 1262 1128 1266 1132
rect 1310 1128 1314 1132
rect 1334 1118 1338 1122
rect 1270 1108 1274 1112
rect 1278 1098 1282 1102
rect 1262 1008 1266 1012
rect 1238 988 1242 992
rect 1254 988 1258 992
rect 1198 958 1202 962
rect 1222 958 1226 962
rect 1318 1088 1322 1092
rect 1342 1078 1346 1082
rect 1294 1068 1298 1072
rect 1326 1068 1330 1072
rect 1278 998 1282 1002
rect 1230 938 1234 942
rect 1270 938 1274 942
rect 1254 918 1258 922
rect 1254 898 1258 902
rect 1302 928 1306 932
rect 1366 1338 1370 1342
rect 1382 1338 1386 1342
rect 1398 1298 1402 1302
rect 1374 1288 1378 1292
rect 1390 1278 1394 1282
rect 1382 1268 1386 1272
rect 1470 1448 1474 1452
rect 1486 1438 1490 1442
rect 1454 1428 1458 1432
rect 1454 1418 1458 1422
rect 1494 1418 1498 1422
rect 1530 1403 1534 1407
rect 1537 1403 1541 1407
rect 1574 1458 1578 1462
rect 1590 1448 1594 1452
rect 1614 1418 1618 1422
rect 1558 1408 1562 1412
rect 1486 1388 1490 1392
rect 1550 1388 1554 1392
rect 1446 1368 1450 1372
rect 1614 1378 1618 1382
rect 1494 1358 1498 1362
rect 1614 1358 1618 1362
rect 1422 1348 1426 1352
rect 1462 1348 1466 1352
rect 1526 1348 1530 1352
rect 1702 1488 1706 1492
rect 1710 1488 1714 1492
rect 1734 1488 1738 1492
rect 1742 1488 1746 1492
rect 1678 1478 1682 1482
rect 1686 1478 1690 1482
rect 1638 1438 1642 1442
rect 1670 1418 1674 1422
rect 1646 1368 1650 1372
rect 1662 1358 1666 1362
rect 1646 1348 1650 1352
rect 1654 1328 1658 1332
rect 1566 1318 1570 1322
rect 1462 1308 1466 1312
rect 1606 1298 1610 1302
rect 1422 1288 1426 1292
rect 1454 1288 1458 1292
rect 1542 1288 1546 1292
rect 1510 1268 1514 1272
rect 1574 1268 1578 1272
rect 1390 1258 1394 1262
rect 1406 1258 1410 1262
rect 1622 1278 1626 1282
rect 1622 1268 1626 1272
rect 1646 1268 1650 1272
rect 1582 1258 1586 1262
rect 1598 1258 1602 1262
rect 1622 1258 1626 1262
rect 1422 1248 1426 1252
rect 1478 1248 1482 1252
rect 1382 1158 1386 1162
rect 1446 1198 1450 1202
rect 1438 1158 1442 1162
rect 1438 1148 1442 1152
rect 1374 1078 1378 1082
rect 1598 1208 1602 1212
rect 1530 1203 1534 1207
rect 1537 1203 1541 1207
rect 1494 1178 1498 1182
rect 1742 1478 1746 1482
rect 1774 1508 1778 1512
rect 1790 1528 1794 1532
rect 1798 1528 1802 1532
rect 1782 1498 1786 1502
rect 1774 1478 1778 1482
rect 1718 1448 1722 1452
rect 1710 1418 1714 1422
rect 1718 1408 1722 1412
rect 1726 1408 1730 1412
rect 1702 1378 1706 1382
rect 1726 1398 1730 1402
rect 1750 1428 1754 1432
rect 1726 1378 1730 1382
rect 1846 1568 1850 1572
rect 1830 1538 1834 1542
rect 1814 1488 1818 1492
rect 1838 1518 1842 1522
rect 1830 1498 1834 1502
rect 1990 1658 1994 1662
rect 1974 1648 1978 1652
rect 1998 1648 2002 1652
rect 2014 1648 2018 1652
rect 1966 1638 1970 1642
rect 1958 1578 1962 1582
rect 1902 1558 1906 1562
rect 1918 1558 1922 1562
rect 1934 1558 1938 1562
rect 1886 1548 1890 1552
rect 1886 1538 1890 1542
rect 1894 1538 1898 1542
rect 1878 1528 1882 1532
rect 1846 1508 1850 1512
rect 1942 1508 1946 1512
rect 1966 1508 1970 1512
rect 1918 1498 1922 1502
rect 1910 1488 1914 1492
rect 1822 1478 1826 1482
rect 1830 1478 1834 1482
rect 1846 1478 1850 1482
rect 1950 1478 1954 1482
rect 1790 1458 1794 1462
rect 1766 1408 1770 1412
rect 1758 1378 1762 1382
rect 1750 1368 1754 1372
rect 1734 1348 1738 1352
rect 1678 1338 1682 1342
rect 1670 1318 1674 1322
rect 1686 1298 1690 1302
rect 1694 1278 1698 1282
rect 1694 1268 1698 1272
rect 1638 1258 1642 1262
rect 1678 1258 1682 1262
rect 1630 1228 1634 1232
rect 1630 1208 1634 1212
rect 1518 1168 1522 1172
rect 1598 1158 1602 1162
rect 1566 1148 1570 1152
rect 1654 1248 1658 1252
rect 1654 1238 1658 1242
rect 1782 1368 1786 1372
rect 1790 1358 1794 1362
rect 1806 1448 1810 1452
rect 1806 1358 1810 1362
rect 1782 1348 1786 1352
rect 1798 1348 1802 1352
rect 1782 1338 1786 1342
rect 1798 1338 1802 1342
rect 1878 1468 1882 1472
rect 1822 1448 1826 1452
rect 1870 1458 1874 1462
rect 1878 1458 1882 1462
rect 1830 1398 1834 1402
rect 1846 1368 1850 1372
rect 1870 1438 1874 1442
rect 1942 1468 1946 1472
rect 1974 1468 1978 1472
rect 1910 1428 1914 1432
rect 1934 1438 1938 1442
rect 1942 1438 1946 1442
rect 1966 1438 1970 1442
rect 1950 1428 1954 1432
rect 1910 1418 1914 1422
rect 1926 1418 1930 1422
rect 1926 1398 1930 1402
rect 2038 1688 2042 1692
rect 2046 1668 2050 1672
rect 2006 1528 2010 1532
rect 1990 1428 1994 1432
rect 1998 1378 2002 1382
rect 1878 1358 1882 1362
rect 1894 1358 1898 1362
rect 1934 1358 1938 1362
rect 1958 1358 1962 1362
rect 1974 1358 1978 1362
rect 1982 1358 1986 1362
rect 1838 1348 1842 1352
rect 1862 1338 1866 1342
rect 1814 1328 1818 1332
rect 1838 1328 1842 1332
rect 1766 1318 1770 1322
rect 1798 1318 1802 1322
rect 1862 1318 1866 1322
rect 1710 1308 1714 1312
rect 1718 1308 1722 1312
rect 1766 1288 1770 1292
rect 1870 1298 1874 1302
rect 1814 1288 1818 1292
rect 1838 1288 1842 1292
rect 1710 1278 1714 1282
rect 1742 1278 1746 1282
rect 1774 1278 1778 1282
rect 1798 1278 1802 1282
rect 1726 1268 1730 1272
rect 1734 1258 1738 1262
rect 1718 1248 1722 1252
rect 1742 1248 1746 1252
rect 1926 1338 1930 1342
rect 1942 1338 1946 1342
rect 1886 1308 1890 1312
rect 1878 1288 1882 1292
rect 1878 1268 1882 1272
rect 2022 1478 2026 1482
rect 2014 1438 2018 1442
rect 2038 1378 2042 1382
rect 2038 1368 2042 1372
rect 1990 1348 1994 1352
rect 2006 1348 2010 1352
rect 1966 1338 1970 1342
rect 1982 1338 1986 1342
rect 2006 1328 2010 1332
rect 1958 1318 1962 1322
rect 1894 1298 1898 1302
rect 1950 1298 1954 1302
rect 1990 1298 1994 1302
rect 1998 1298 2002 1302
rect 2030 1298 2034 1302
rect 1902 1288 1906 1292
rect 1934 1278 1938 1282
rect 2030 1278 2034 1282
rect 1958 1268 1962 1272
rect 2014 1268 2018 1272
rect 2038 1268 2042 1272
rect 1918 1258 1922 1262
rect 1942 1258 1946 1262
rect 1822 1248 1826 1252
rect 1854 1248 1858 1252
rect 1742 1238 1746 1242
rect 1790 1238 1794 1242
rect 1854 1238 1858 1242
rect 1702 1188 1706 1192
rect 1670 1178 1674 1182
rect 1694 1168 1698 1172
rect 1630 1158 1634 1162
rect 1646 1158 1650 1162
rect 1662 1158 1666 1162
rect 1646 1148 1650 1152
rect 1574 1138 1578 1142
rect 1606 1138 1610 1142
rect 1622 1138 1626 1142
rect 1558 1128 1562 1132
rect 1654 1128 1658 1132
rect 1358 1068 1362 1072
rect 1366 1068 1370 1072
rect 1454 1068 1458 1072
rect 1374 1058 1378 1062
rect 1334 1048 1338 1052
rect 1350 1048 1354 1052
rect 1326 1018 1330 1022
rect 1326 928 1330 932
rect 1342 918 1346 922
rect 1302 898 1306 902
rect 1318 898 1322 902
rect 1334 898 1338 902
rect 1222 868 1226 872
rect 1254 868 1258 872
rect 1142 858 1146 862
rect 1190 858 1194 862
rect 1318 868 1322 872
rect 1398 1038 1402 1042
rect 1366 1018 1370 1022
rect 1446 988 1450 992
rect 1486 988 1490 992
rect 1502 988 1506 992
rect 1382 948 1386 952
rect 1398 948 1402 952
rect 1414 948 1418 952
rect 1382 938 1386 942
rect 1406 918 1410 922
rect 1374 908 1378 912
rect 1350 888 1354 892
rect 1286 858 1290 862
rect 1166 848 1170 852
rect 1158 828 1162 832
rect 1150 788 1154 792
rect 1158 788 1162 792
rect 1182 778 1186 782
rect 1134 758 1138 762
rect 1070 738 1074 742
rect 1126 738 1130 742
rect 1022 728 1026 732
rect 1018 703 1022 707
rect 1025 703 1029 707
rect 1022 658 1026 662
rect 1014 578 1018 582
rect 1166 748 1170 752
rect 1198 768 1202 772
rect 1334 828 1338 832
rect 1310 768 1314 772
rect 1246 747 1250 751
rect 1302 748 1306 752
rect 1246 738 1250 742
rect 1094 728 1098 732
rect 1134 728 1138 732
rect 1150 728 1154 732
rect 1158 728 1162 732
rect 1062 698 1066 702
rect 1182 688 1186 692
rect 1198 678 1202 682
rect 1230 668 1234 672
rect 1110 658 1114 662
rect 1046 648 1050 652
rect 1038 628 1042 632
rect 1030 568 1034 572
rect 958 458 962 462
rect 974 458 978 462
rect 934 448 938 452
rect 982 438 986 442
rect 894 428 898 432
rect 894 398 898 402
rect 870 388 874 392
rect 854 368 858 372
rect 838 338 842 342
rect 782 318 786 322
rect 806 318 810 322
rect 822 318 826 322
rect 774 298 778 302
rect 766 268 770 272
rect 798 268 802 272
rect 774 238 778 242
rect 782 218 786 222
rect 798 208 802 212
rect 726 138 730 142
rect 686 108 690 112
rect 798 148 802 152
rect 742 128 746 132
rect 686 78 690 82
rect 702 78 706 82
rect 790 128 794 132
rect 758 98 762 102
rect 830 298 834 302
rect 822 288 826 292
rect 830 278 834 282
rect 990 368 994 372
rect 974 348 978 352
rect 870 338 874 342
rect 934 338 938 342
rect 1030 528 1034 532
rect 1038 528 1042 532
rect 1018 503 1022 507
rect 1025 503 1029 507
rect 1126 648 1130 652
rect 1070 618 1074 622
rect 1150 608 1154 612
rect 1102 558 1106 562
rect 1118 548 1122 552
rect 1134 548 1138 552
rect 1286 728 1290 732
rect 1262 668 1266 672
rect 1294 668 1298 672
rect 1438 938 1442 942
rect 1454 938 1458 942
rect 1470 938 1474 942
rect 1582 1118 1586 1122
rect 1590 1118 1594 1122
rect 1638 1118 1642 1122
rect 1558 1098 1562 1102
rect 1622 1098 1626 1102
rect 1598 1088 1602 1092
rect 1646 1078 1650 1082
rect 1606 1068 1610 1072
rect 1638 1068 1642 1072
rect 1606 1058 1610 1062
rect 1654 1058 1658 1062
rect 1542 1028 1546 1032
rect 1606 1028 1610 1032
rect 1530 1003 1534 1007
rect 1537 1003 1541 1007
rect 1518 978 1522 982
rect 1494 938 1498 942
rect 1510 938 1514 942
rect 1614 968 1618 972
rect 1630 958 1634 962
rect 1662 958 1666 962
rect 1566 948 1570 952
rect 1526 938 1530 942
rect 1438 928 1442 932
rect 1478 928 1482 932
rect 1470 898 1474 902
rect 1366 878 1370 882
rect 1422 878 1426 882
rect 1326 758 1330 762
rect 1350 758 1354 762
rect 1358 758 1362 762
rect 1350 728 1354 732
rect 1326 678 1330 682
rect 1342 678 1346 682
rect 1246 648 1250 652
rect 1166 578 1170 582
rect 1190 558 1194 562
rect 1166 548 1170 552
rect 1278 618 1282 622
rect 1438 868 1442 872
rect 1510 928 1514 932
rect 1550 928 1554 932
rect 1502 908 1506 912
rect 1502 888 1506 892
rect 1518 888 1522 892
rect 1598 928 1602 932
rect 1606 928 1610 932
rect 1614 918 1618 922
rect 1758 1158 1762 1162
rect 1758 1138 1762 1142
rect 1678 1088 1682 1092
rect 1710 1088 1714 1092
rect 1734 1088 1738 1092
rect 1694 1078 1698 1082
rect 1750 1078 1754 1082
rect 1766 1078 1770 1082
rect 1702 1058 1706 1062
rect 1710 1058 1714 1062
rect 1726 1058 1730 1062
rect 1694 998 1698 1002
rect 1678 978 1682 982
rect 1694 958 1698 962
rect 1670 948 1674 952
rect 1662 938 1666 942
rect 1886 1208 1890 1212
rect 1910 1208 1914 1212
rect 1838 1188 1842 1192
rect 1886 1138 1890 1142
rect 1910 1138 1914 1142
rect 1854 1098 1858 1102
rect 1870 1068 1874 1072
rect 1806 1048 1810 1052
rect 1838 1048 1842 1052
rect 1718 958 1722 962
rect 1710 938 1714 942
rect 1678 928 1682 932
rect 1582 898 1586 902
rect 1638 898 1642 902
rect 1454 858 1458 862
rect 1494 858 1498 862
rect 1518 858 1522 862
rect 1478 848 1482 852
rect 1470 838 1474 842
rect 1374 768 1378 772
rect 1398 768 1402 772
rect 1414 768 1418 772
rect 1446 738 1450 742
rect 1398 728 1402 732
rect 1430 728 1434 732
rect 1366 718 1370 722
rect 1398 698 1402 702
rect 1414 698 1418 702
rect 1406 688 1410 692
rect 1366 668 1370 672
rect 1310 658 1314 662
rect 1326 658 1330 662
rect 1358 658 1362 662
rect 1374 658 1378 662
rect 1318 648 1322 652
rect 1302 558 1306 562
rect 1294 548 1298 552
rect 1158 538 1162 542
rect 1238 538 1242 542
rect 1294 538 1298 542
rect 1318 538 1322 542
rect 1078 528 1082 532
rect 1126 528 1130 532
rect 1054 518 1058 522
rect 1102 518 1106 522
rect 1078 498 1082 502
rect 1086 498 1090 502
rect 1150 508 1154 512
rect 1110 498 1114 502
rect 1094 488 1098 492
rect 1038 468 1042 472
rect 1046 468 1050 472
rect 1030 448 1034 452
rect 1038 438 1042 442
rect 1006 368 1010 372
rect 1142 488 1146 492
rect 1078 468 1082 472
rect 1126 468 1130 472
rect 1166 528 1170 532
rect 1174 528 1178 532
rect 1174 508 1178 512
rect 1222 508 1226 512
rect 1174 498 1178 502
rect 1278 468 1282 472
rect 1054 458 1058 462
rect 1070 458 1074 462
rect 1126 458 1130 462
rect 1054 428 1058 432
rect 998 338 1002 342
rect 1054 338 1058 342
rect 990 328 994 332
rect 990 318 994 322
rect 1006 318 1010 322
rect 1038 318 1042 322
rect 1054 318 1058 322
rect 1062 318 1066 322
rect 854 278 858 282
rect 870 278 874 282
rect 878 278 882 282
rect 950 278 954 282
rect 846 268 850 272
rect 862 268 866 272
rect 830 258 834 262
rect 814 228 818 232
rect 814 198 818 202
rect 910 268 914 272
rect 942 268 946 272
rect 966 268 970 272
rect 974 268 978 272
rect 982 268 986 272
rect 886 258 890 262
rect 894 258 898 262
rect 934 258 938 262
rect 878 248 882 252
rect 870 218 874 222
rect 862 158 866 162
rect 822 138 826 142
rect 782 78 786 82
rect 806 78 810 82
rect 838 98 842 102
rect 846 68 850 72
rect 878 158 882 162
rect 902 248 906 252
rect 942 218 946 222
rect 894 208 898 212
rect 942 208 946 212
rect 1018 303 1022 307
rect 1025 303 1029 307
rect 1006 258 1010 262
rect 1006 208 1010 212
rect 958 188 962 192
rect 1022 178 1026 182
rect 1006 168 1010 172
rect 998 148 1002 152
rect 982 138 986 142
rect 990 128 994 132
rect 910 98 914 102
rect 878 88 882 92
rect 1018 103 1022 107
rect 1025 103 1029 107
rect 1046 268 1050 272
rect 1134 448 1138 452
rect 1142 448 1146 452
rect 1262 448 1266 452
rect 1110 398 1114 402
rect 1094 368 1098 372
rect 1118 368 1122 372
rect 1110 348 1114 352
rect 1102 338 1106 342
rect 1134 338 1138 342
rect 1278 438 1282 442
rect 1222 428 1226 432
rect 1206 368 1210 372
rect 1150 338 1154 342
rect 1158 328 1162 332
rect 1126 318 1130 322
rect 1118 308 1122 312
rect 1078 288 1082 292
rect 1046 228 1050 232
rect 1062 228 1066 232
rect 1030 88 1034 92
rect 1038 88 1042 92
rect 1118 278 1122 282
rect 1190 298 1194 302
rect 1214 278 1218 282
rect 1094 268 1098 272
rect 1134 268 1138 272
rect 1166 268 1170 272
rect 1134 258 1138 262
rect 1126 248 1130 252
rect 1246 398 1250 402
rect 1294 518 1298 522
rect 1334 648 1338 652
rect 1350 618 1354 622
rect 1334 548 1338 552
rect 1374 648 1378 652
rect 1366 588 1370 592
rect 1366 558 1370 562
rect 1334 528 1338 532
rect 1326 508 1330 512
rect 1350 488 1354 492
rect 1334 478 1338 482
rect 1454 678 1458 682
rect 1462 678 1466 682
rect 1446 668 1450 672
rect 1534 828 1538 832
rect 1530 803 1534 807
rect 1537 803 1541 807
rect 1486 788 1490 792
rect 1534 788 1538 792
rect 1502 768 1506 772
rect 1478 758 1482 762
rect 1494 758 1498 762
rect 1550 738 1554 742
rect 1590 888 1594 892
rect 1646 888 1650 892
rect 1654 878 1658 882
rect 1646 868 1650 872
rect 1566 858 1570 862
rect 1590 848 1594 852
rect 1630 808 1634 812
rect 1566 768 1570 772
rect 1574 758 1578 762
rect 1590 758 1594 762
rect 1606 758 1610 762
rect 1582 738 1586 742
rect 1598 738 1602 742
rect 1606 738 1610 742
rect 1542 728 1546 732
rect 1542 688 1546 692
rect 1478 678 1482 682
rect 1502 668 1506 672
rect 1518 668 1522 672
rect 1534 668 1538 672
rect 1510 658 1514 662
rect 1614 688 1618 692
rect 1606 678 1610 682
rect 1582 668 1586 672
rect 1478 648 1482 652
rect 1414 598 1418 602
rect 1530 603 1534 607
rect 1537 603 1541 607
rect 1534 588 1538 592
rect 1398 548 1402 552
rect 1510 548 1514 552
rect 1390 538 1394 542
rect 1422 538 1426 542
rect 1590 548 1594 552
rect 1438 528 1442 532
rect 1590 518 1594 522
rect 1598 508 1602 512
rect 1438 488 1442 492
rect 1454 488 1458 492
rect 1518 488 1522 492
rect 1478 478 1482 482
rect 1502 478 1506 482
rect 1558 478 1562 482
rect 1406 468 1410 472
rect 1454 468 1458 472
rect 1486 468 1490 472
rect 1598 468 1602 472
rect 1302 458 1306 462
rect 1382 458 1386 462
rect 1286 388 1290 392
rect 1286 348 1290 352
rect 1302 348 1306 352
rect 1278 338 1282 342
rect 1254 268 1258 272
rect 1302 318 1306 322
rect 1462 458 1466 462
rect 1398 398 1402 402
rect 1326 388 1330 392
rect 1350 368 1354 372
rect 1366 368 1370 372
rect 1358 358 1362 362
rect 1334 338 1338 342
rect 1422 338 1426 342
rect 1430 328 1434 332
rect 1366 318 1370 322
rect 1278 268 1282 272
rect 1334 268 1338 272
rect 1422 308 1426 312
rect 1446 278 1450 282
rect 1486 448 1490 452
rect 1558 448 1562 452
rect 1510 438 1514 442
rect 1486 428 1490 432
rect 1530 403 1534 407
rect 1537 403 1541 407
rect 1542 388 1546 392
rect 1510 298 1514 302
rect 1462 268 1466 272
rect 1478 268 1482 272
rect 1206 258 1210 262
rect 1246 258 1250 262
rect 1270 258 1274 262
rect 1318 258 1322 262
rect 1406 258 1410 262
rect 1446 258 1450 262
rect 1206 248 1210 252
rect 1246 248 1250 252
rect 1182 228 1186 232
rect 1190 228 1194 232
rect 1302 238 1306 242
rect 1158 208 1162 212
rect 1294 208 1298 212
rect 1150 168 1154 172
rect 1150 158 1154 162
rect 1174 158 1178 162
rect 1222 158 1226 162
rect 1158 148 1162 152
rect 1190 148 1194 152
rect 1182 138 1186 142
rect 1254 138 1258 142
rect 1142 128 1146 132
rect 1102 118 1106 122
rect 1206 118 1210 122
rect 1078 78 1082 82
rect 1366 158 1370 162
rect 1358 148 1362 152
rect 1118 88 1122 92
rect 1190 88 1194 92
rect 1222 88 1226 92
rect 1310 88 1314 92
rect 1334 88 1338 92
rect 1374 88 1378 92
rect 1166 78 1170 82
rect 1214 78 1218 82
rect 1310 78 1314 82
rect 918 68 922 72
rect 942 68 946 72
rect 1054 68 1058 72
rect 1086 68 1090 72
rect 1174 68 1178 72
rect 1374 68 1378 72
rect 438 58 442 62
rect 470 58 474 62
rect 582 58 586 62
rect 654 58 658 62
rect 862 58 866 62
rect 958 58 962 62
rect 1566 438 1570 442
rect 1638 648 1642 652
rect 1630 638 1634 642
rect 1662 858 1666 862
rect 1718 918 1722 922
rect 1710 858 1714 862
rect 1710 848 1714 852
rect 1822 1038 1826 1042
rect 1806 958 1810 962
rect 1998 1258 2002 1262
rect 1982 1238 1986 1242
rect 2046 1238 2050 1242
rect 2022 1158 2026 1162
rect 1990 1148 1994 1152
rect 1982 1118 1986 1122
rect 1966 1108 1970 1112
rect 1926 1078 1930 1082
rect 2014 1098 2018 1102
rect 1974 1068 1978 1072
rect 1998 1068 2002 1072
rect 1910 1058 1914 1062
rect 1950 1058 1954 1062
rect 1878 1038 1882 1042
rect 1902 1028 1906 1032
rect 1902 1008 1906 1012
rect 1822 948 1826 952
rect 1750 938 1754 942
rect 1734 928 1738 932
rect 1742 898 1746 902
rect 1782 918 1786 922
rect 1774 908 1778 912
rect 1782 898 1786 902
rect 1758 888 1762 892
rect 1766 888 1770 892
rect 1790 888 1794 892
rect 1790 878 1794 882
rect 1774 858 1778 862
rect 1710 838 1714 842
rect 1726 838 1730 842
rect 1678 778 1682 782
rect 1726 768 1730 772
rect 1654 758 1658 762
rect 1678 758 1682 762
rect 1758 768 1762 772
rect 1894 938 1898 942
rect 1910 868 1914 872
rect 1846 858 1850 862
rect 1854 848 1858 852
rect 1814 758 1818 762
rect 1766 748 1770 752
rect 1798 748 1802 752
rect 1734 738 1738 742
rect 1790 738 1794 742
rect 1694 728 1698 732
rect 1686 718 1690 722
rect 1654 668 1658 672
rect 1662 668 1666 672
rect 1654 638 1658 642
rect 1814 708 1818 712
rect 1846 708 1850 712
rect 1806 698 1810 702
rect 1822 698 1826 702
rect 1694 668 1698 672
rect 1950 1048 1954 1052
rect 1926 918 1930 922
rect 2046 1048 2050 1052
rect 2022 1028 2026 1032
rect 2022 1018 2026 1022
rect 2006 958 2010 962
rect 1982 938 1986 942
rect 1966 878 1970 882
rect 1926 868 1930 872
rect 1950 858 1954 862
rect 1918 848 1922 852
rect 1934 848 1938 852
rect 1910 838 1914 842
rect 1902 828 1906 832
rect 1958 748 1962 752
rect 1862 738 1866 742
rect 1918 738 1922 742
rect 1942 738 1946 742
rect 1870 698 1874 702
rect 1878 688 1882 692
rect 1862 668 1866 672
rect 1910 668 1914 672
rect 1678 658 1682 662
rect 1734 658 1738 662
rect 1822 658 1826 662
rect 1926 658 1930 662
rect 1686 648 1690 652
rect 1670 588 1674 592
rect 1694 558 1698 562
rect 1758 648 1762 652
rect 1774 648 1778 652
rect 1750 638 1754 642
rect 1766 618 1770 622
rect 1846 638 1850 642
rect 1742 548 1746 552
rect 1614 488 1618 492
rect 1646 458 1650 462
rect 1646 438 1650 442
rect 1622 398 1626 402
rect 1606 388 1610 392
rect 1630 388 1634 392
rect 1590 378 1594 382
rect 1622 378 1626 382
rect 1558 358 1562 362
rect 1422 178 1426 182
rect 1462 178 1466 182
rect 1414 168 1418 172
rect 1530 203 1534 207
rect 1537 203 1541 207
rect 1462 168 1466 172
rect 1614 308 1618 312
rect 1574 298 1578 302
rect 1702 538 1706 542
rect 1662 528 1666 532
rect 1710 528 1714 532
rect 1750 528 1754 532
rect 1670 508 1674 512
rect 1742 508 1746 512
rect 1702 498 1706 502
rect 1670 488 1674 492
rect 1678 478 1682 482
rect 1654 428 1658 432
rect 1726 488 1730 492
rect 1798 548 1802 552
rect 1790 538 1794 542
rect 1846 538 1850 542
rect 1886 648 1890 652
rect 1918 648 1922 652
rect 1910 638 1914 642
rect 1894 618 1898 622
rect 1926 628 1930 632
rect 1926 558 1930 562
rect 1862 548 1866 552
rect 1902 548 1906 552
rect 1782 478 1786 482
rect 1886 478 1890 482
rect 1958 728 1962 732
rect 2006 858 2010 862
rect 1998 748 2002 752
rect 2038 828 2042 832
rect 1998 738 2002 742
rect 1990 728 1994 732
rect 1974 698 1978 702
rect 1950 678 1954 682
rect 1966 678 1970 682
rect 1990 678 1994 682
rect 1966 668 1970 672
rect 1958 658 1962 662
rect 1950 618 1954 622
rect 2006 688 2010 692
rect 2014 678 2018 682
rect 2030 668 2034 672
rect 2022 658 2026 662
rect 2006 558 2010 562
rect 1926 548 1930 552
rect 1942 548 1946 552
rect 1966 548 1970 552
rect 2038 548 2042 552
rect 1926 538 1930 542
rect 1918 498 1922 502
rect 1902 468 1906 472
rect 1774 458 1778 462
rect 1846 458 1850 462
rect 1878 458 1882 462
rect 1678 448 1682 452
rect 1678 418 1682 422
rect 1702 418 1706 422
rect 1742 418 1746 422
rect 1734 408 1738 412
rect 1678 398 1682 402
rect 1670 388 1674 392
rect 1694 378 1698 382
rect 1718 378 1722 382
rect 1694 348 1698 352
rect 1734 368 1738 372
rect 1742 358 1746 362
rect 1782 358 1786 362
rect 1918 428 1922 432
rect 1846 418 1850 422
rect 1862 418 1866 422
rect 1918 418 1922 422
rect 1814 368 1818 372
rect 1838 368 1842 372
rect 1774 348 1778 352
rect 1806 348 1810 352
rect 1694 338 1698 342
rect 1662 328 1666 332
rect 1598 278 1602 282
rect 1630 278 1634 282
rect 1670 278 1674 282
rect 1678 278 1682 282
rect 1558 268 1562 272
rect 1606 268 1610 272
rect 1566 258 1570 262
rect 1646 258 1650 262
rect 1558 168 1562 172
rect 1438 148 1442 152
rect 1550 148 1554 152
rect 1430 138 1434 142
rect 1462 138 1466 142
rect 1446 118 1450 122
rect 1622 248 1626 252
rect 1638 248 1642 252
rect 1678 248 1682 252
rect 1638 188 1642 192
rect 1598 178 1602 182
rect 1622 178 1626 182
rect 1630 168 1634 172
rect 1598 138 1602 142
rect 1654 158 1658 162
rect 1726 318 1730 322
rect 1686 168 1690 172
rect 1790 338 1794 342
rect 1766 318 1770 322
rect 1790 288 1794 292
rect 1894 358 1898 362
rect 1846 328 1850 332
rect 1814 318 1818 322
rect 1806 268 1810 272
rect 1814 268 1818 272
rect 1758 258 1762 262
rect 1782 178 1786 182
rect 1806 178 1810 182
rect 1694 148 1698 152
rect 1734 148 1738 152
rect 1654 138 1658 142
rect 1678 138 1682 142
rect 1510 128 1514 132
rect 1630 128 1634 132
rect 1622 98 1626 102
rect 1534 88 1538 92
rect 1566 88 1570 92
rect 1590 88 1594 92
rect 1614 88 1618 92
rect 1606 78 1610 82
rect 1134 58 1138 62
rect 1166 58 1170 62
rect 1214 58 1218 62
rect 1734 108 1738 112
rect 1822 228 1826 232
rect 1886 338 1890 342
rect 1870 298 1874 302
rect 1990 528 1994 532
rect 1950 478 1954 482
rect 2006 518 2010 522
rect 2030 528 2034 532
rect 2014 508 2018 512
rect 2014 498 2018 502
rect 2022 478 2026 482
rect 2030 468 2034 472
rect 2006 458 2010 462
rect 2014 458 2018 462
rect 2038 458 2042 462
rect 1958 388 1962 392
rect 1942 368 1946 372
rect 1878 278 1882 282
rect 1926 278 1930 282
rect 1902 268 1906 272
rect 1926 258 1930 262
rect 1942 248 1946 252
rect 1974 308 1978 312
rect 1958 218 1962 222
rect 1950 188 1954 192
rect 1854 168 1858 172
rect 1870 168 1874 172
rect 1830 148 1834 152
rect 1862 148 1866 152
rect 1766 108 1770 112
rect 1718 78 1722 82
rect 1766 68 1770 72
rect 1862 118 1866 122
rect 1870 118 1874 122
rect 1862 68 1866 72
rect 1966 178 1970 182
rect 1982 268 1986 272
rect 1990 218 1994 222
rect 1998 198 2002 202
rect 2014 328 2018 332
rect 2030 258 2034 262
rect 1990 98 1994 102
rect 1982 88 1986 92
rect 2014 98 2018 102
rect 486 48 490 52
rect 662 48 666 52
rect 678 48 682 52
rect 782 48 786 52
rect 1126 48 1130 52
rect 1158 48 1162 52
rect 1206 48 1210 52
rect 1270 48 1274 52
rect 414 38 418 42
rect 2022 88 2026 92
rect 2022 58 2026 62
rect 1990 8 1994 12
rect 2014 8 2018 12
rect 498 3 502 7
rect 505 3 509 7
rect 1530 3 1534 7
rect 1537 3 1541 7
<< metal3 >>
rect 496 1803 498 1807
rect 502 1803 505 1807
rect 510 1803 512 1807
rect 1528 1803 1530 1807
rect 1534 1803 1537 1807
rect 1542 1803 1544 1807
rect -26 1798 -22 1802
rect 10 1798 174 1801
rect 818 1798 830 1801
rect -26 1791 -23 1798
rect -26 1788 14 1791
rect 26 1788 33 1791
rect 58 1788 118 1791
rect 122 1788 918 1791
rect 30 1782 33 1788
rect -26 1781 -22 1782
rect -26 1778 6 1781
rect 1950 1768 1966 1771
rect 2078 1771 2082 1772
rect 2010 1768 2082 1771
rect 1950 1762 1953 1768
rect -26 1761 -22 1762
rect -26 1758 126 1761
rect 1934 1752 1937 1758
rect 14 1748 150 1751
rect 610 1748 670 1751
rect 922 1748 1214 1751
rect 1218 1748 1665 1751
rect 2078 1751 2082 1752
rect 2050 1748 2082 1751
rect -26 1741 -22 1742
rect 14 1741 17 1748
rect -26 1738 17 1741
rect 354 1738 374 1741
rect 658 1738 774 1741
rect 798 1741 801 1748
rect 1662 1742 1665 1748
rect 798 1738 854 1741
rect 914 1738 942 1741
rect 1146 1738 1350 1741
rect 1466 1738 1486 1741
rect 1490 1738 1510 1741
rect 1666 1738 1670 1741
rect 534 1728 662 1731
rect 1006 1731 1009 1738
rect 930 1728 1150 1731
rect 1218 1728 1230 1731
rect 1234 1728 1294 1731
rect 1390 1731 1393 1738
rect 1390 1728 1438 1731
rect 1442 1728 1510 1731
rect 1574 1731 1577 1738
rect 1514 1728 1734 1731
rect 1822 1731 1825 1738
rect 1738 1728 1825 1731
rect 1950 1731 1953 1738
rect 1938 1728 1953 1731
rect 2018 1728 2022 1731
rect -26 1721 -22 1722
rect 406 1721 409 1728
rect 534 1722 537 1728
rect 1966 1722 1969 1728
rect -26 1718 409 1721
rect 450 1718 534 1721
rect 690 1718 710 1721
rect 826 1718 1118 1721
rect 1194 1718 1222 1721
rect 1902 1712 1905 1718
rect 498 1708 510 1711
rect 578 1708 822 1711
rect 1962 1708 2006 1711
rect 1016 1703 1018 1707
rect 1022 1703 1025 1707
rect 1030 1703 1032 1707
rect 146 1698 190 1701
rect 306 1698 486 1701
rect 1266 1698 1406 1701
rect 170 1688 358 1691
rect 978 1688 990 1691
rect 1618 1688 1670 1691
rect 1810 1688 1846 1691
rect 94 1681 97 1688
rect 94 1678 110 1681
rect 114 1678 286 1681
rect 994 1678 1006 1681
rect 1010 1678 1062 1681
rect 1066 1678 1094 1681
rect 1250 1678 1254 1681
rect 1258 1678 1342 1681
rect 1902 1681 1905 1688
rect 1882 1678 1905 1681
rect 2038 1681 2041 1688
rect 1986 1678 2041 1681
rect 402 1668 574 1671
rect 818 1668 902 1671
rect 1050 1668 1070 1671
rect 1162 1668 1174 1671
rect 1178 1668 1246 1671
rect 1258 1668 1286 1671
rect 1542 1668 1550 1671
rect 1842 1668 1902 1671
rect 1906 1668 1910 1671
rect 1914 1668 2046 1671
rect 1542 1662 1545 1668
rect 170 1658 230 1661
rect 522 1658 534 1661
rect 650 1658 678 1661
rect 682 1658 1110 1661
rect 1114 1658 1126 1661
rect 1146 1658 1182 1661
rect 1210 1658 1286 1661
rect 1594 1658 1614 1661
rect 1898 1658 1990 1661
rect 2014 1652 2017 1658
rect 354 1648 582 1651
rect 586 1648 662 1651
rect 666 1648 790 1651
rect 946 1648 1065 1651
rect 982 1642 985 1648
rect 1062 1642 1065 1648
rect 1086 1648 1118 1651
rect 1218 1648 1254 1651
rect 1802 1648 1838 1651
rect 1842 1648 1870 1651
rect 1978 1648 1998 1651
rect 1086 1642 1089 1648
rect 290 1638 718 1641
rect 1178 1638 1206 1641
rect 1330 1638 1454 1641
rect 1650 1638 1654 1641
rect 1658 1638 1966 1641
rect 1970 1638 1974 1641
rect 466 1628 734 1631
rect 1074 1628 1166 1631
rect 250 1618 590 1621
rect 594 1618 614 1621
rect 618 1618 710 1621
rect 762 1618 798 1621
rect 802 1618 822 1621
rect 1030 1618 1150 1621
rect 1030 1612 1033 1618
rect 1230 1612 1233 1618
rect 754 1608 782 1611
rect 496 1603 498 1607
rect 502 1603 505 1607
rect 510 1603 512 1607
rect 1528 1603 1530 1607
rect 1534 1603 1537 1607
rect 1542 1603 1544 1607
rect 554 1598 774 1601
rect 1698 1598 1718 1601
rect 34 1588 54 1591
rect 842 1588 846 1591
rect 1218 1588 1246 1591
rect 630 1582 633 1588
rect 1130 1578 1166 1581
rect 1170 1578 1278 1581
rect 1738 1578 1958 1581
rect -26 1571 -22 1572
rect 6 1571 9 1578
rect -26 1568 9 1571
rect 614 1568 758 1571
rect 974 1571 977 1578
rect 778 1568 977 1571
rect 1090 1568 1142 1571
rect 1154 1568 1174 1571
rect 50 1558 214 1561
rect 526 1561 529 1568
rect 614 1562 617 1568
rect 442 1558 529 1561
rect 578 1558 614 1561
rect 714 1558 742 1561
rect 746 1558 1158 1561
rect 1194 1558 1294 1561
rect 1846 1561 1849 1568
rect 1794 1558 1849 1561
rect 1922 1558 1934 1561
rect -26 1551 -22 1552
rect -26 1548 30 1551
rect 42 1548 174 1551
rect 218 1548 526 1551
rect 530 1548 566 1551
rect 630 1551 633 1558
rect 602 1548 633 1551
rect 1066 1548 1070 1551
rect 1122 1548 1126 1551
rect 1586 1548 1622 1551
rect 1810 1548 1886 1551
rect 1902 1551 1905 1558
rect 1890 1548 1905 1551
rect 450 1538 590 1541
rect 594 1538 646 1541
rect 846 1541 849 1548
rect 778 1538 849 1541
rect 962 1538 1006 1541
rect 1010 1538 1046 1541
rect 1154 1538 1214 1541
rect 1338 1538 1510 1541
rect 1514 1538 1518 1541
rect 1834 1538 1886 1541
rect 1898 1538 1902 1541
rect 138 1528 142 1531
rect 146 1528 166 1531
rect 170 1528 358 1531
rect 362 1528 382 1531
rect 1102 1531 1105 1538
rect 386 1528 1105 1531
rect 1134 1531 1137 1538
rect 1134 1528 1382 1531
rect 1386 1528 1470 1531
rect 1694 1531 1697 1538
rect 1694 1528 1734 1531
rect 1738 1528 1750 1531
rect 1794 1528 1798 1531
rect 1882 1528 2006 1531
rect 602 1518 654 1521
rect 1098 1518 1110 1521
rect 1114 1518 1190 1521
rect 1234 1518 1361 1521
rect 1442 1518 1462 1521
rect 1682 1518 1838 1521
rect 1358 1512 1361 1518
rect 114 1508 614 1511
rect 674 1508 694 1511
rect 1074 1508 1198 1511
rect 1202 1508 1238 1511
rect 1290 1508 1334 1511
rect 1778 1508 1846 1511
rect 1946 1508 1966 1511
rect 750 1502 753 1508
rect 1016 1503 1018 1507
rect 1022 1503 1025 1507
rect 1030 1503 1032 1507
rect 154 1498 390 1501
rect 562 1498 718 1501
rect 1122 1498 1246 1501
rect 1250 1498 1254 1501
rect 1354 1498 1406 1501
rect 1602 1498 1630 1501
rect 1634 1498 1782 1501
rect 1826 1498 1830 1501
rect 1842 1498 1918 1501
rect 106 1488 142 1491
rect 282 1488 622 1491
rect 866 1488 950 1491
rect 1258 1488 1430 1491
rect 1530 1488 1542 1491
rect 1698 1488 1702 1491
rect 1714 1488 1734 1491
rect 1746 1488 1814 1491
rect 1818 1488 1910 1491
rect 630 1482 633 1488
rect 98 1478 166 1481
rect 170 1478 254 1481
rect 266 1478 358 1481
rect 498 1478 542 1481
rect 546 1478 550 1481
rect 758 1481 761 1488
rect 666 1478 761 1481
rect 842 1478 846 1481
rect 1194 1478 1206 1481
rect 1218 1478 1310 1481
rect 1466 1478 1518 1481
rect 1522 1478 1614 1481
rect 1618 1478 1678 1481
rect 1690 1478 1742 1481
rect 1834 1478 1846 1481
rect 1954 1478 2022 1481
rect 42 1468 110 1471
rect 114 1468 121 1471
rect 130 1468 174 1471
rect 194 1468 246 1471
rect 358 1471 361 1478
rect 358 1468 446 1471
rect 466 1468 558 1471
rect 578 1468 582 1471
rect 642 1468 862 1471
rect 898 1468 958 1471
rect 1050 1468 1118 1471
rect 1186 1468 1238 1471
rect 1378 1468 1742 1471
rect 1774 1471 1777 1478
rect 1822 1471 1825 1478
rect 1774 1468 1801 1471
rect 1822 1468 1878 1471
rect 1882 1468 1942 1471
rect 1946 1468 1974 1471
rect 122 1458 142 1461
rect 146 1458 182 1461
rect 186 1458 246 1461
rect 522 1458 542 1461
rect 1002 1458 1038 1461
rect 1066 1458 1222 1461
rect 1226 1458 1273 1461
rect 1298 1458 1318 1461
rect 1322 1458 1366 1461
rect 1370 1458 1438 1461
rect 1442 1458 1550 1461
rect 1554 1458 1574 1461
rect 1578 1458 1790 1461
rect 1798 1461 1801 1468
rect 1798 1458 1854 1461
rect 1874 1458 1878 1461
rect 1270 1452 1273 1458
rect 130 1448 134 1451
rect 138 1448 214 1451
rect 522 1448 542 1451
rect 602 1448 1022 1451
rect 1026 1448 1054 1451
rect 1154 1448 1174 1451
rect 1210 1448 1254 1451
rect 1282 1448 1294 1451
rect 1474 1448 1590 1451
rect 1714 1448 1718 1451
rect 1826 1448 1830 1451
rect 1834 1448 1902 1451
rect 1906 1448 1937 1451
rect 106 1438 134 1441
rect 194 1438 206 1441
rect 594 1438 1102 1441
rect 1178 1438 1206 1441
rect 1234 1438 1262 1441
rect 1266 1438 1286 1441
rect 1354 1438 1422 1441
rect 1490 1438 1638 1441
rect 1806 1441 1809 1448
rect 1934 1442 1937 1448
rect 2014 1442 2017 1448
rect 1642 1438 1809 1441
rect 1858 1438 1870 1441
rect 1946 1438 1966 1441
rect 226 1428 558 1431
rect 562 1428 582 1431
rect 586 1428 870 1431
rect 874 1428 894 1431
rect 898 1428 1006 1431
rect 1010 1428 1070 1431
rect 1186 1428 1230 1431
rect 1234 1428 1246 1431
rect 1250 1428 1270 1431
rect 1282 1428 1454 1431
rect 1458 1428 1750 1431
rect 1914 1428 1950 1431
rect 1994 1428 1998 1431
rect 202 1418 302 1421
rect 1162 1418 1382 1421
rect 1386 1418 1454 1421
rect 1498 1418 1614 1421
rect 1674 1418 1710 1421
rect 1714 1418 1910 1421
rect 1930 1418 1958 1421
rect 678 1412 681 1418
rect 930 1408 1182 1411
rect 1234 1408 1286 1411
rect 1314 1408 1470 1411
rect 1562 1408 1718 1411
rect 1730 1408 1734 1411
rect 1770 1408 1998 1411
rect 496 1403 498 1407
rect 502 1403 505 1407
rect 510 1403 512 1407
rect 1528 1403 1530 1407
rect 1534 1403 1537 1407
rect 1542 1403 1544 1407
rect 786 1398 806 1401
rect 810 1398 1038 1401
rect 1042 1398 1078 1401
rect 1082 1398 1158 1401
rect 1162 1398 1414 1401
rect 1730 1398 1734 1401
rect 1834 1398 1926 1401
rect 210 1388 214 1391
rect 1082 1388 1094 1391
rect 1102 1388 1278 1391
rect 1290 1388 1486 1391
rect 1554 1388 1761 1391
rect 706 1378 1038 1381
rect 1102 1381 1105 1388
rect 1758 1382 1761 1388
rect 1058 1378 1105 1381
rect 1114 1378 1134 1381
rect 1138 1378 1278 1381
rect 1282 1378 1406 1381
rect 1618 1378 1702 1381
rect 1706 1378 1726 1381
rect 1766 1378 1998 1381
rect 2026 1378 2038 1381
rect 466 1368 526 1371
rect 1018 1368 1190 1371
rect 1266 1368 1270 1371
rect 1450 1368 1646 1371
rect 1766 1371 1769 1378
rect 1754 1368 1769 1371
rect 1786 1368 1846 1371
rect 2034 1368 2038 1371
rect 918 1362 921 1368
rect 1254 1362 1257 1368
rect 138 1358 382 1361
rect 690 1358 734 1361
rect 962 1358 1022 1361
rect 1026 1358 1206 1361
rect 1322 1358 1342 1361
rect 1486 1358 1494 1361
rect 1498 1358 1614 1361
rect 1794 1358 1806 1361
rect 1882 1358 1894 1361
rect 1898 1358 1934 1361
rect 1962 1358 1974 1361
rect 1986 1358 1990 1361
rect 186 1348 190 1351
rect 426 1348 470 1351
rect 474 1348 494 1351
rect 654 1351 657 1358
rect 570 1348 657 1351
rect 662 1352 665 1358
rect 706 1348 742 1351
rect 778 1348 790 1351
rect 886 1351 889 1358
rect 886 1348 942 1351
rect 1098 1348 1142 1351
rect 1218 1348 1230 1351
rect 1314 1348 1358 1351
rect 1378 1348 1382 1351
rect 1426 1348 1462 1351
rect 1662 1351 1665 1358
rect 1650 1348 1665 1351
rect 1738 1348 1782 1351
rect 1786 1348 1793 1351
rect 1802 1348 1838 1351
rect 1842 1348 1977 1351
rect 1994 1348 2006 1351
rect 162 1338 254 1341
rect 394 1338 414 1341
rect 530 1338 638 1341
rect 642 1338 662 1341
rect 666 1338 694 1341
rect 698 1338 710 1341
rect 714 1338 934 1341
rect 938 1338 974 1341
rect 978 1338 1286 1341
rect 1370 1338 1382 1341
rect 1526 1341 1529 1348
rect 1974 1342 1977 1348
rect 1522 1338 1529 1341
rect 1682 1338 1782 1341
rect 1786 1338 1790 1341
rect 1802 1338 1862 1341
rect 1930 1338 1942 1341
rect 1946 1338 1966 1341
rect 1978 1338 1982 1341
rect 94 1331 97 1338
rect 34 1328 230 1331
rect 234 1328 297 1331
rect 410 1328 422 1331
rect 478 1331 481 1338
rect 458 1328 481 1331
rect 562 1328 806 1331
rect 810 1328 985 1331
rect 1258 1328 1318 1331
rect 1346 1328 1654 1331
rect 1818 1328 1838 1331
rect 1842 1328 2006 1331
rect 294 1322 297 1328
rect 982 1322 985 1328
rect 402 1318 446 1321
rect 530 1318 598 1321
rect 674 1318 678 1321
rect 682 1318 758 1321
rect 762 1318 806 1321
rect 818 1318 822 1321
rect 1002 1318 1078 1321
rect 1106 1318 1358 1321
rect 1570 1318 1670 1321
rect 1770 1318 1798 1321
rect 1866 1318 1958 1321
rect 114 1308 414 1311
rect 434 1308 438 1311
rect 450 1308 558 1311
rect 762 1308 766 1311
rect 786 1308 870 1311
rect 874 1308 926 1311
rect 1050 1308 1150 1311
rect 1162 1308 1174 1311
rect 1178 1308 1350 1311
rect 1466 1308 1710 1311
rect 1722 1308 1886 1311
rect 2078 1311 2082 1312
rect 1890 1308 2082 1311
rect 1016 1303 1018 1307
rect 1022 1303 1025 1307
rect 1030 1303 1032 1307
rect 154 1298 446 1301
rect 826 1298 870 1301
rect 874 1298 918 1301
rect 1154 1298 1182 1301
rect 1402 1298 1606 1301
rect 1610 1298 1686 1301
rect 1690 1298 1870 1301
rect 1898 1298 1950 1301
rect 1954 1298 1966 1301
rect 1986 1298 1990 1301
rect 2002 1298 2030 1301
rect 274 1288 294 1291
rect 298 1288 390 1291
rect 394 1288 430 1291
rect 442 1288 454 1291
rect 458 1288 465 1291
rect 494 1291 497 1298
rect 490 1288 497 1291
rect 506 1288 574 1291
rect 706 1288 894 1291
rect 906 1288 990 1291
rect 1378 1288 1422 1291
rect 1458 1288 1542 1291
rect 1562 1288 1697 1291
rect 1762 1288 1766 1291
rect 1818 1288 1822 1291
rect 1842 1288 1878 1291
rect 1898 1288 1902 1291
rect 1906 1288 2046 1291
rect 110 1281 113 1288
rect 1094 1282 1097 1288
rect 1158 1282 1161 1288
rect 1694 1282 1697 1288
rect 110 1278 150 1281
rect 202 1278 286 1281
rect 314 1278 406 1281
rect 442 1278 470 1281
rect 506 1278 598 1281
rect 610 1278 678 1281
rect 834 1278 838 1281
rect 850 1278 854 1281
rect 874 1278 886 1281
rect 1314 1278 1390 1281
rect 1626 1278 1649 1281
rect 1714 1278 1742 1281
rect 1778 1278 1798 1281
rect 1838 1281 1841 1288
rect 1802 1278 1841 1281
rect 1870 1278 1934 1281
rect 2026 1278 2030 1281
rect 58 1268 118 1271
rect 258 1268 310 1271
rect 314 1268 425 1271
rect 474 1268 478 1271
rect 490 1268 577 1271
rect 586 1268 590 1271
rect 666 1268 670 1271
rect 706 1268 862 1271
rect 866 1268 1038 1271
rect 1042 1268 1046 1271
rect 1066 1268 1078 1271
rect 1086 1271 1089 1278
rect 1646 1272 1649 1278
rect 1086 1268 1102 1271
rect 1386 1268 1390 1271
rect 1514 1268 1574 1271
rect 1594 1268 1622 1271
rect 1690 1268 1694 1271
rect 1870 1271 1873 1278
rect 1730 1268 1873 1271
rect 1882 1268 1958 1271
rect 2018 1268 2038 1271
rect 2078 1271 2082 1272
rect 2050 1268 2082 1271
rect 130 1258 134 1261
rect 158 1258 214 1261
rect 250 1258 262 1261
rect 266 1258 342 1261
rect 346 1258 350 1261
rect 370 1258 406 1261
rect 422 1261 425 1268
rect 422 1258 510 1261
rect 574 1261 577 1268
rect 574 1258 662 1261
rect 710 1258 766 1261
rect 810 1258 862 1261
rect 946 1258 998 1261
rect 1010 1258 1054 1261
rect 1058 1258 1110 1261
rect 1130 1258 1230 1261
rect 1394 1258 1398 1261
rect 1402 1258 1406 1261
rect 1586 1258 1598 1261
rect 1618 1258 1622 1261
rect 1642 1258 1678 1261
rect 1682 1258 1734 1261
rect 1746 1258 1918 1261
rect 1934 1258 1942 1261
rect 1946 1258 1998 1261
rect 158 1252 161 1258
rect 710 1252 713 1258
rect 202 1248 278 1251
rect 378 1248 542 1251
rect 546 1248 678 1251
rect 762 1248 830 1251
rect 1082 1248 1310 1251
rect 1354 1248 1422 1251
rect 1426 1248 1478 1251
rect 1658 1248 1718 1251
rect 1746 1248 1822 1251
rect 1826 1248 1838 1251
rect 2078 1251 2082 1252
rect 1858 1248 2082 1251
rect 374 1242 377 1248
rect 1718 1242 1721 1248
rect 442 1238 462 1241
rect 538 1238 558 1241
rect 562 1238 654 1241
rect 658 1238 742 1241
rect 746 1238 846 1241
rect 866 1238 1134 1241
rect 1170 1238 1222 1241
rect 1658 1238 1710 1241
rect 1730 1238 1742 1241
rect 1794 1238 1854 1241
rect 1986 1238 2046 1241
rect 450 1228 478 1231
rect 498 1228 534 1231
rect 550 1228 630 1231
rect 682 1228 782 1231
rect 794 1228 1062 1231
rect 1106 1228 1174 1231
rect 550 1222 553 1228
rect 1630 1222 1633 1228
rect 442 1218 470 1221
rect 754 1218 766 1221
rect 1122 1218 1230 1221
rect 1886 1212 1889 1218
rect 1910 1212 1913 1218
rect 690 1208 814 1211
rect 1634 1208 1734 1211
rect 496 1203 498 1207
rect 502 1203 505 1207
rect 510 1203 512 1207
rect 1528 1203 1530 1207
rect 1534 1203 1537 1207
rect 1542 1203 1544 1207
rect 1598 1202 1601 1208
rect 1242 1198 1446 1201
rect 618 1188 638 1191
rect 842 1188 1078 1191
rect 1090 1188 1702 1191
rect 402 1178 462 1181
rect 586 1178 638 1181
rect 642 1178 646 1181
rect 858 1178 862 1181
rect 874 1178 1297 1181
rect 1498 1178 1625 1181
rect 1838 1181 1841 1188
rect 1674 1178 1841 1181
rect 1294 1172 1297 1178
rect 434 1168 582 1171
rect 586 1168 918 1171
rect 1330 1168 1518 1171
rect 1622 1171 1625 1178
rect 1622 1168 1694 1171
rect 226 1158 422 1161
rect 538 1158 654 1161
rect 658 1158 862 1161
rect 918 1161 921 1168
rect 1190 1162 1193 1168
rect 882 1158 926 1161
rect 970 1158 1062 1161
rect 1194 1158 1206 1161
rect 1442 1158 1454 1161
rect 1518 1161 1521 1168
rect 1518 1158 1574 1161
rect 1578 1158 1598 1161
rect 1602 1158 1630 1161
rect 1650 1158 1662 1161
rect 1762 1158 2022 1161
rect 222 1151 225 1158
rect 210 1148 225 1151
rect 306 1148 382 1151
rect 418 1148 422 1151
rect 442 1148 649 1151
rect 770 1148 798 1151
rect 866 1148 958 1151
rect 962 1148 998 1151
rect 1094 1151 1097 1158
rect 1382 1152 1385 1158
rect 1058 1148 1097 1151
rect 1298 1148 1302 1151
rect 1514 1148 1566 1151
rect 1570 1148 1606 1151
rect 1910 1148 1990 1151
rect 110 1141 113 1148
rect 270 1141 273 1148
rect 34 1138 273 1141
rect 426 1138 470 1141
rect 490 1138 518 1141
rect 522 1138 542 1141
rect 546 1138 558 1141
rect 610 1138 638 1141
rect 646 1141 649 1148
rect 646 1138 894 1141
rect 1058 1138 1078 1141
rect 1082 1138 1110 1141
rect 1178 1138 1182 1141
rect 1258 1138 1294 1141
rect 1314 1138 1318 1141
rect 1438 1141 1441 1148
rect 1646 1142 1649 1148
rect 1910 1142 1913 1148
rect 1438 1138 1569 1141
rect 1578 1138 1606 1141
rect 1610 1138 1622 1141
rect 1762 1138 1886 1141
rect 146 1128 230 1131
rect 378 1128 406 1131
rect 410 1128 478 1131
rect 530 1128 614 1131
rect 642 1128 678 1131
rect 682 1128 766 1131
rect 978 1128 1022 1131
rect 1162 1128 1262 1131
rect 1314 1128 1462 1131
rect 1566 1131 1569 1138
rect 1566 1128 1593 1131
rect 1642 1128 1654 1131
rect 1758 1131 1761 1138
rect 1754 1128 1761 1131
rect 614 1121 617 1128
rect 614 1118 654 1121
rect 658 1118 678 1121
rect 826 1118 1126 1121
rect 1154 1118 1206 1121
rect 1210 1118 1334 1121
rect 1558 1121 1561 1128
rect 1590 1122 1593 1128
rect 1558 1118 1582 1121
rect 1642 1118 1942 1121
rect 1946 1118 1982 1121
rect 458 1108 486 1111
rect 554 1108 702 1111
rect 1250 1108 1270 1111
rect 1290 1108 1966 1111
rect 1016 1103 1018 1107
rect 1022 1103 1025 1107
rect 1030 1103 1032 1107
rect 170 1098 398 1101
rect 474 1098 550 1101
rect 554 1098 582 1101
rect 650 1098 670 1101
rect 714 1098 718 1101
rect 730 1098 822 1101
rect 1242 1098 1278 1101
rect 1282 1098 1510 1101
rect 1562 1098 1622 1101
rect 1858 1098 1934 1101
rect 1938 1098 2014 1101
rect 58 1088 182 1091
rect 278 1088 358 1091
rect 418 1088 574 1091
rect 706 1088 830 1091
rect 858 1088 878 1091
rect 882 1088 902 1091
rect 1218 1088 1318 1091
rect 1730 1088 1734 1091
rect 10 1078 174 1081
rect 222 1081 225 1088
rect 278 1082 281 1088
rect 646 1082 649 1088
rect 178 1078 225 1081
rect 258 1078 262 1081
rect 314 1078 318 1081
rect 402 1078 406 1081
rect 418 1078 438 1081
rect 466 1078 470 1081
rect 690 1078 694 1081
rect 722 1078 726 1081
rect 802 1078 886 1081
rect 942 1081 945 1088
rect 906 1078 945 1081
rect 1298 1078 1342 1081
rect 1346 1078 1374 1081
rect 1598 1081 1601 1088
rect 1598 1078 1646 1081
rect 1678 1081 1681 1088
rect 1666 1078 1681 1081
rect 1698 1078 1702 1081
rect 1710 1081 1713 1088
rect 1710 1078 1750 1081
rect 1770 1078 1926 1081
rect 130 1068 174 1071
rect 250 1068 302 1071
rect 306 1068 350 1071
rect 354 1068 374 1071
rect 378 1068 422 1071
rect 426 1068 454 1071
rect 514 1068 542 1071
rect 674 1068 750 1071
rect 870 1068 894 1071
rect 930 1068 934 1071
rect 1002 1068 1046 1071
rect 1134 1071 1137 1078
rect 1134 1068 1206 1071
rect 1298 1068 1326 1071
rect 1330 1068 1358 1071
rect 1370 1068 1454 1071
rect 1474 1068 1606 1071
rect 1610 1068 1638 1071
rect 1658 1068 1870 1071
rect 1978 1068 1998 1071
rect 574 1062 577 1068
rect 870 1062 873 1068
rect 138 1058 150 1061
rect 274 1058 321 1061
rect 330 1058 414 1061
rect 522 1058 526 1061
rect 690 1058 694 1061
rect 730 1058 854 1061
rect 962 1058 966 1061
rect 970 1058 1022 1061
rect 1030 1058 1102 1061
rect 1242 1058 1337 1061
rect 1378 1058 1606 1061
rect 1658 1058 1702 1061
rect 1706 1058 1710 1061
rect 1722 1058 1726 1061
rect 1914 1058 1926 1061
rect 1930 1058 1950 1061
rect 318 1052 321 1058
rect 422 1052 425 1058
rect 430 1052 433 1058
rect 1030 1052 1033 1058
rect 1334 1052 1337 1058
rect 74 1048 129 1051
rect 126 1042 129 1048
rect 682 1048 694 1051
rect 914 1048 974 1051
rect 1338 1048 1350 1051
rect 1802 1048 1806 1051
rect 1842 1048 1950 1051
rect 2042 1048 2046 1051
rect 2078 1051 2082 1052
rect 2050 1048 2082 1051
rect 214 1042 217 1048
rect 854 1042 857 1048
rect 274 1038 334 1041
rect 402 1038 438 1041
rect 570 1038 694 1041
rect 906 1038 918 1041
rect 986 1038 1046 1041
rect 1130 1038 1214 1041
rect 1218 1038 1398 1041
rect 1826 1038 1878 1041
rect 110 1031 113 1038
rect 110 1028 206 1031
rect 210 1028 374 1031
rect 562 1028 910 1031
rect 1138 1028 1142 1031
rect 1170 1028 1174 1031
rect 1178 1028 1542 1031
rect 1610 1028 1902 1031
rect 2010 1028 2022 1031
rect 586 1018 734 1021
rect 1330 1018 1366 1021
rect 1490 1018 2022 1021
rect 806 1012 809 1018
rect 610 1008 758 1011
rect 810 1008 894 1011
rect 1026 1008 1262 1011
rect 1906 1008 1910 1011
rect 496 1003 498 1007
rect 502 1003 505 1007
rect 510 1003 512 1007
rect 1528 1003 1530 1007
rect 1534 1003 1537 1007
rect 1542 1003 1544 1007
rect 650 998 718 1001
rect 722 998 766 1001
rect 1158 998 1278 1001
rect 622 992 625 998
rect 10 988 30 991
rect 282 988 382 991
rect 410 988 478 991
rect 722 988 782 991
rect 874 988 934 991
rect 1158 991 1161 998
rect 1694 992 1697 998
rect 938 988 1161 991
rect 1242 988 1254 991
rect 1258 988 1446 991
rect 1450 988 1486 991
rect 1490 988 1502 991
rect 302 978 478 981
rect 814 981 817 988
rect 762 978 817 981
rect 922 978 926 981
rect 994 978 1150 981
rect 1238 981 1241 988
rect 1170 978 1241 981
rect 1522 978 1678 981
rect 302 972 305 978
rect 742 972 745 978
rect 862 972 865 978
rect 498 968 534 971
rect 538 968 582 971
rect 658 968 726 971
rect 770 968 790 971
rect 794 968 830 971
rect 1082 968 1182 971
rect 1266 968 1614 971
rect 1626 968 1721 971
rect 186 958 222 961
rect 226 958 230 961
rect 366 961 369 968
rect 1718 962 1721 968
rect 366 958 398 961
rect 418 958 454 961
rect 474 958 1198 961
rect 1202 958 1222 961
rect 1226 958 1630 961
rect 1634 958 1662 961
rect 1798 958 1806 961
rect 1810 958 2006 961
rect 130 948 198 951
rect 338 948 545 951
rect 554 948 646 951
rect 650 948 662 951
rect 738 948 745 951
rect 794 948 830 951
rect 858 948 934 951
rect 938 948 966 951
rect 1058 948 1086 951
rect 1138 948 1158 951
rect 1162 948 1174 951
rect 1386 948 1390 951
rect 1402 948 1414 951
rect 1466 948 1566 951
rect 1570 948 1670 951
rect 1694 951 1697 958
rect 1694 948 1822 951
rect 206 941 209 948
rect 318 941 321 948
rect 162 938 321 941
rect 458 938 462 941
rect 482 938 486 941
rect 542 941 545 948
rect 742 942 745 948
rect 1454 942 1457 948
rect 542 938 574 941
rect 594 938 598 941
rect 642 938 646 941
rect 786 938 798 941
rect 826 938 990 941
rect 1002 938 1126 941
rect 1130 938 1230 941
rect 1274 938 1305 941
rect 1386 938 1438 941
rect 1474 938 1494 941
rect 1506 938 1510 941
rect 1606 938 1622 941
rect 1658 938 1662 941
rect 1714 938 1750 941
rect 1898 938 1982 941
rect 274 928 286 931
rect 334 931 337 938
rect 334 928 358 931
rect 402 928 406 931
rect 534 931 537 938
rect 1302 932 1305 938
rect 426 928 537 931
rect 762 928 838 931
rect 850 928 854 931
rect 898 928 902 931
rect 914 928 1158 931
rect 1330 928 1409 931
rect 1442 928 1478 931
rect 1526 931 1529 938
rect 1606 932 1609 938
rect 1514 928 1529 931
rect 1546 928 1550 931
rect 1594 928 1598 931
rect 1682 928 1734 931
rect 1406 922 1409 928
rect 210 918 310 921
rect 314 918 422 921
rect 450 918 598 921
rect 650 918 686 921
rect 738 918 806 921
rect 810 918 1158 921
rect 1258 918 1342 921
rect 1414 918 1614 921
rect 1722 918 1782 921
rect 1786 918 1926 921
rect 218 908 278 911
rect 298 908 374 911
rect 378 908 558 911
rect 618 908 670 911
rect 730 908 758 911
rect 858 908 886 911
rect 1050 908 1374 911
rect 1414 911 1417 918
rect 1378 908 1417 911
rect 1506 908 1598 911
rect 1602 908 1774 911
rect 1016 903 1018 907
rect 1022 903 1025 907
rect 1030 903 1032 907
rect 154 898 198 901
rect 306 898 310 901
rect 314 898 342 901
rect 346 898 374 901
rect 378 898 430 901
rect 434 898 662 901
rect 826 898 870 901
rect 1038 898 1254 901
rect 1306 898 1318 901
rect 1322 898 1334 901
rect 1474 898 1582 901
rect 1642 898 1742 901
rect 1746 898 1782 901
rect 154 888 174 891
rect 258 888 326 891
rect 442 888 454 891
rect 506 888 590 891
rect 610 888 638 891
rect 642 888 654 891
rect 658 888 702 891
rect 722 888 742 891
rect 834 888 838 891
rect 850 888 854 891
rect 1038 891 1041 898
rect 906 888 1041 891
rect 1050 888 1054 891
rect 1154 888 1158 891
rect 1354 888 1478 891
rect 1482 888 1502 891
rect 1522 888 1590 891
rect 1602 888 1646 891
rect 1762 888 1766 891
rect 1770 888 1790 891
rect 10 878 102 881
rect 106 878 182 881
rect 194 878 230 881
rect 374 881 377 888
rect 282 878 377 881
rect 442 878 625 881
rect 634 878 654 881
rect 658 878 1006 881
rect 1042 878 1366 881
rect 1426 878 1654 881
rect 1794 878 1966 881
rect 254 871 257 878
rect 90 868 257 871
rect 362 868 390 871
rect 394 868 446 871
rect 622 871 625 878
rect 622 868 750 871
rect 834 868 878 871
rect 930 868 990 871
rect 1142 868 1222 871
rect 1258 868 1318 871
rect 1454 868 1646 871
rect 1706 868 1713 871
rect 1790 871 1793 878
rect 1770 868 1793 871
rect 70 861 73 868
rect 70 858 118 861
rect 130 858 134 861
rect 138 858 158 861
rect 178 858 222 861
rect 346 858 401 861
rect 410 858 454 861
rect 554 859 606 861
rect 550 858 606 859
rect 746 858 750 861
rect 778 858 782 861
rect 798 861 801 868
rect 990 862 993 868
rect 1062 862 1065 868
rect 1142 862 1145 868
rect 1438 862 1441 868
rect 1454 862 1457 868
rect 1710 862 1713 868
rect 1910 862 1913 868
rect 798 858 822 861
rect 842 858 870 861
rect 1010 858 1038 861
rect 1194 858 1286 861
rect 1498 858 1518 861
rect 1570 858 1662 861
rect 1778 858 1846 861
rect 1926 861 1929 868
rect 1926 858 1950 861
rect 2010 858 2014 861
rect 398 852 401 858
rect 1006 852 1009 858
rect 618 848 630 851
rect 690 848 718 851
rect 722 848 785 851
rect 794 848 806 851
rect 1034 848 1102 851
rect 1170 848 1478 851
rect 1594 848 1622 851
rect 1666 848 1710 851
rect 1714 848 1721 851
rect 1858 848 1918 851
rect 1922 848 1934 851
rect 782 842 785 848
rect 394 838 606 841
rect 866 838 910 841
rect 914 838 966 841
rect 970 838 1470 841
rect 1474 838 1590 841
rect 1594 838 1710 841
rect 1730 838 1910 841
rect 162 828 182 831
rect 186 828 582 831
rect 626 828 646 831
rect 726 831 729 838
rect 658 828 729 831
rect 834 828 1158 831
rect 1338 828 1534 831
rect 1538 828 1686 831
rect 1690 828 1902 831
rect 1906 828 2038 831
rect 98 818 414 821
rect 530 818 582 821
rect 618 818 918 821
rect 946 818 950 821
rect 1630 812 1633 818
rect 122 808 134 811
rect 138 808 142 811
rect 146 808 182 811
rect 186 808 470 811
rect 706 808 726 811
rect 834 808 942 811
rect 496 803 498 807
rect 502 803 505 807
rect 510 803 512 807
rect 1528 803 1530 807
rect 1534 803 1537 807
rect 1542 803 1544 807
rect 242 798 310 801
rect 426 798 478 801
rect 962 798 974 801
rect 226 788 270 791
rect 458 788 502 791
rect 770 788 774 791
rect 810 788 1150 791
rect 1162 788 1190 791
rect 1490 788 1534 791
rect 426 778 526 781
rect 534 781 537 788
rect 534 778 614 781
rect 698 778 862 781
rect 866 778 998 781
rect 1002 778 1006 781
rect 1010 778 1182 781
rect 1194 778 1678 781
rect 306 768 398 771
rect 402 768 526 771
rect 730 768 838 771
rect 922 768 934 771
rect 962 768 990 771
rect 1202 768 1310 771
rect 1378 768 1398 771
rect 1402 768 1406 771
rect 1418 768 1502 771
rect 1506 768 1566 771
rect 1610 768 1726 771
rect 1762 768 1817 771
rect 450 758 470 761
rect 490 758 494 761
rect 514 758 542 761
rect 550 761 553 768
rect 1814 762 1817 768
rect 546 758 553 761
rect 682 758 702 761
rect 714 758 718 761
rect 754 758 878 761
rect 890 758 974 761
rect 1050 758 1070 761
rect 1074 758 1086 761
rect 1090 758 1118 761
rect 1138 758 1150 761
rect 1330 758 1350 761
rect 1362 758 1478 761
rect 1498 758 1574 761
rect 1586 758 1590 761
rect 1610 758 1614 761
rect 1658 758 1678 761
rect 58 748 134 751
rect 214 751 217 758
rect 470 752 473 758
rect 170 748 217 751
rect 370 748 438 751
rect 482 748 510 751
rect 514 748 550 751
rect 610 748 625 751
rect 142 742 145 748
rect 122 738 142 741
rect 146 738 182 741
rect 334 741 337 748
rect 590 742 593 748
rect 622 742 625 748
rect 666 748 670 751
rect 730 748 734 751
rect 746 748 750 751
rect 762 748 766 751
rect 794 748 846 751
rect 890 748 934 751
rect 970 748 1054 751
rect 1066 748 1166 751
rect 250 738 337 741
rect 466 738 534 741
rect 630 741 633 748
rect 1250 748 1294 751
rect 1306 748 1598 751
rect 1602 748 1766 751
rect 1770 748 1798 751
rect 1962 748 1998 751
rect 1942 742 1945 748
rect 630 738 662 741
rect 674 738 678 741
rect 714 738 734 741
rect 754 738 761 741
rect 778 738 782 741
rect 826 738 830 741
rect 842 738 894 741
rect 914 738 918 741
rect 978 738 1070 741
rect 1130 738 1238 741
rect 1250 738 1433 741
rect 1442 738 1446 741
rect 1546 738 1550 741
rect 1574 738 1582 741
rect 1586 738 1598 741
rect 1610 738 1702 741
rect 1706 738 1734 741
rect 1794 738 1862 741
rect 1946 738 1998 741
rect 758 732 761 738
rect 1430 732 1433 738
rect 178 728 182 731
rect 318 728 350 731
rect 442 728 478 731
rect 678 728 686 731
rect 690 728 718 731
rect 786 728 798 731
rect 810 728 830 731
rect 850 728 950 731
rect 1026 728 1094 731
rect 1114 728 1134 731
rect 1154 728 1158 731
rect 1162 728 1286 731
rect 1298 728 1350 731
rect 1390 728 1398 731
rect 1402 728 1422 731
rect 1450 728 1542 731
rect 1546 728 1553 731
rect 1642 728 1694 731
rect 1918 731 1921 738
rect 1918 728 1934 731
rect 1962 728 1990 731
rect 318 722 321 728
rect 330 718 606 721
rect 610 718 694 721
rect 858 718 886 721
rect 906 718 1166 721
rect 1170 718 1222 721
rect 1370 718 1686 721
rect 1690 718 1806 721
rect 154 708 286 711
rect 522 708 878 711
rect 1818 708 1846 711
rect 1016 703 1018 707
rect 1022 703 1025 707
rect 1030 703 1032 707
rect 250 698 286 701
rect 466 698 566 701
rect 586 698 721 701
rect 762 698 790 701
rect 1066 698 1398 701
rect 1418 698 1510 701
rect 1810 698 1822 701
rect 1874 698 1974 701
rect 106 688 150 691
rect 154 688 486 691
rect 578 688 590 691
rect 658 688 710 691
rect 718 691 721 698
rect 718 688 758 691
rect 762 688 870 691
rect 986 688 990 691
rect 1546 688 1614 691
rect 1950 688 2006 691
rect 194 678 270 681
rect 282 678 294 681
rect 466 678 478 681
rect 482 678 489 681
rect 506 678 553 681
rect 594 678 646 681
rect 694 678 702 681
rect 706 678 726 681
rect 1182 681 1185 688
rect 874 678 1185 681
rect 1194 678 1198 681
rect 1230 678 1326 681
rect 1346 678 1350 681
rect 1406 681 1409 688
rect 1406 678 1454 681
rect 1466 678 1470 681
rect 1482 678 1606 681
rect 1878 681 1881 688
rect 1682 678 1881 681
rect 1950 682 1953 688
rect 2014 682 2017 691
rect 1970 678 1990 681
rect 106 668 142 671
rect 266 668 302 671
rect 334 671 337 678
rect 550 672 553 678
rect 1230 672 1233 678
rect 334 668 422 671
rect 426 668 470 671
rect 490 668 510 671
rect 522 668 526 671
rect 642 668 702 671
rect 706 668 750 671
rect 850 668 854 671
rect 930 668 934 671
rect 994 668 998 671
rect 1266 668 1286 671
rect 1298 668 1366 671
rect 1450 668 1494 671
rect 1498 668 1502 671
rect 1522 668 1526 671
rect 1538 668 1582 671
rect 1666 668 1694 671
rect 1866 668 1910 671
rect 1914 668 1966 671
rect 1970 668 2030 671
rect 58 658 118 661
rect 138 658 142 661
rect 146 658 150 661
rect 186 658 254 661
rect 290 658 302 661
rect 330 658 374 661
rect 466 658 542 661
rect 706 658 710 661
rect 818 658 902 661
rect 938 658 1022 661
rect 1114 658 1310 661
rect 1330 658 1358 661
rect 1378 658 1510 661
rect 1514 658 1614 661
rect 1654 661 1657 668
rect 1650 658 1657 661
rect 1682 658 1686 661
rect 1738 658 1822 661
rect 1826 658 1921 661
rect 1930 658 1934 661
rect 1954 658 1958 661
rect 2018 658 2022 661
rect 566 652 569 658
rect 1918 652 1921 658
rect 66 648 166 651
rect 290 648 326 651
rect 554 648 558 651
rect 738 648 838 651
rect 962 648 966 651
rect 1050 648 1126 651
rect 1130 648 1246 651
rect 1274 648 1318 651
rect 1322 648 1334 651
rect 1338 648 1374 651
rect 1482 648 1638 651
rect 1690 648 1758 651
rect 1778 648 1886 651
rect 314 638 326 641
rect 414 638 422 641
rect 426 638 462 641
rect 526 641 529 648
rect 526 638 582 641
rect 774 638 846 641
rect 866 638 886 641
rect 938 638 1630 641
rect 1658 638 1750 641
rect 1850 638 1910 641
rect 774 632 777 638
rect 418 628 742 631
rect 858 628 1038 631
rect 1242 628 1926 631
rect 306 618 649 621
rect 666 618 838 621
rect 882 618 902 621
rect 1074 618 1262 621
rect 1282 618 1350 621
rect 1362 618 1766 621
rect 1898 618 1950 621
rect 98 608 446 611
rect 602 608 622 611
rect 646 611 649 618
rect 646 608 886 611
rect 890 608 1150 611
rect 1154 608 1390 611
rect 496 603 498 607
rect 502 603 505 607
rect 510 603 512 607
rect 1528 603 1530 607
rect 1534 603 1537 607
rect 1542 603 1544 607
rect 794 598 870 601
rect 986 598 1414 601
rect 130 588 262 591
rect 266 588 382 591
rect 434 588 606 591
rect 610 588 686 591
rect 1042 588 1182 591
rect 1186 588 1366 591
rect 1370 588 1486 591
rect 1538 588 1670 591
rect 250 578 414 581
rect 474 578 574 581
rect 578 578 630 581
rect 770 578 790 581
rect 794 578 814 581
rect 1018 578 1166 581
rect 1166 572 1169 578
rect 146 568 214 571
rect 346 568 350 571
rect 474 568 566 571
rect 634 568 830 571
rect 834 568 846 571
rect 1034 568 1102 571
rect 582 562 585 568
rect 2006 562 2009 568
rect 186 558 198 561
rect 202 558 222 561
rect 346 558 374 561
rect 378 558 398 561
rect 410 558 510 561
rect 562 558 582 561
rect 586 558 878 561
rect 882 558 894 561
rect 898 558 910 561
rect 930 558 966 561
rect 1106 558 1190 561
rect 1306 558 1366 561
rect 1650 558 1694 561
rect 1930 558 2006 561
rect 194 548 246 551
rect 306 548 374 551
rect 530 548 590 551
rect 594 548 598 551
rect 622 548 657 551
rect 714 548 766 551
rect 778 548 798 551
rect 802 548 1118 551
rect 1122 548 1134 551
rect 1170 548 1190 551
rect 1194 548 1294 551
rect 1402 548 1510 551
rect 1594 548 1705 551
rect 1746 548 1798 551
rect 1802 548 1862 551
rect 1890 548 1902 551
rect 1906 548 1926 551
rect 1946 548 1966 551
rect 1970 548 2038 551
rect 2078 548 2082 552
rect 622 542 625 548
rect 654 542 657 548
rect 34 538 113 541
rect 138 538 198 541
rect 394 538 598 541
rect 634 538 638 541
rect 754 538 1118 541
rect 1122 538 1158 541
rect 1178 538 1238 541
rect 1298 538 1318 541
rect 1334 541 1337 548
rect 1702 542 1705 548
rect 1334 538 1390 541
rect 1394 538 1422 541
rect 1794 538 1846 541
rect 1930 538 1934 541
rect 2078 541 2081 548
rect 1938 538 2081 541
rect 110 532 113 538
rect 570 528 678 531
rect 706 528 766 531
rect 830 528 870 531
rect 882 528 902 531
rect 938 528 998 531
rect 1002 528 1030 531
rect 1042 528 1078 531
rect 1170 528 1174 531
rect 1338 528 1438 531
rect 1442 528 1638 531
rect 1666 528 1710 531
rect 1754 528 1990 531
rect 2026 528 2030 531
rect 830 522 833 528
rect 82 518 86 521
rect 842 518 1046 521
rect 1058 518 1102 521
rect 1126 521 1129 528
rect 1126 518 1174 521
rect 1298 518 1590 521
rect 2010 518 2038 521
rect 42 508 110 511
rect 130 508 390 511
rect 578 508 590 511
rect 602 508 838 511
rect 850 508 886 511
rect 890 508 918 511
rect 1146 508 1150 511
rect 1178 508 1222 511
rect 1330 508 1598 511
rect 1674 508 1742 511
rect 2018 508 2046 511
rect 1016 503 1018 507
rect 1022 503 1025 507
rect 1030 503 1032 507
rect 1086 502 1089 508
rect 730 498 870 501
rect 906 498 958 501
rect 1050 498 1078 501
rect 1114 498 1174 501
rect 1706 498 1918 501
rect 1930 498 2014 501
rect 242 488 326 491
rect 330 488 518 491
rect 538 488 606 491
rect 874 488 878 491
rect 914 488 918 491
rect 942 488 950 491
rect 954 488 1094 491
rect 1146 488 1350 491
rect 1354 488 1438 491
rect 1458 488 1518 491
rect 1522 488 1614 491
rect 1618 488 1670 491
rect 1730 488 2038 491
rect 226 478 318 481
rect 322 478 350 481
rect 394 478 646 481
rect 754 478 822 481
rect 834 478 1334 481
rect 1490 478 1502 481
rect 1562 478 1678 481
rect 1786 478 1886 481
rect 1954 478 2014 481
rect 2018 478 2022 481
rect 454 472 457 478
rect 1478 472 1481 478
rect 18 468 30 471
rect 98 468 126 471
rect 378 468 422 471
rect 498 468 774 471
rect 850 468 926 471
rect 954 468 1038 471
rect 1050 468 1054 471
rect 1066 468 1078 471
rect 1090 468 1126 471
rect 1138 468 1278 471
rect 1458 468 1478 471
rect 1490 468 1550 471
rect 1602 468 1902 471
rect 2026 468 2030 471
rect 2078 471 2082 472
rect 2042 468 2082 471
rect 122 458 126 461
rect 154 458 166 461
rect 226 459 278 461
rect 226 458 281 459
rect 354 458 374 461
rect 450 458 614 461
rect 618 458 710 461
rect 806 461 809 468
rect 846 461 849 468
rect 806 458 849 461
rect 962 458 966 461
rect 978 458 982 461
rect 1010 458 1054 461
rect 1074 458 1126 461
rect 1130 458 1166 461
rect 1170 458 1302 461
rect 1306 458 1382 461
rect 1406 461 1409 468
rect 1406 458 1462 461
rect 1498 458 1646 461
rect 1650 458 1774 461
rect 1850 458 1878 461
rect 1962 458 2006 461
rect 2018 458 2038 461
rect 862 452 865 458
rect 186 448 230 451
rect 234 448 494 451
rect 530 448 550 451
rect 554 448 822 451
rect 898 448 934 451
rect 1002 448 1030 451
rect 1138 448 1142 451
rect 1146 448 1158 451
rect 1266 448 1270 451
rect 1490 448 1494 451
rect 1562 448 1646 451
rect 2078 451 2082 452
rect 1682 448 2082 451
rect 1278 442 1281 448
rect 194 438 222 441
rect 522 438 534 441
rect 754 438 982 441
rect 1042 438 1086 441
rect 1514 438 1566 441
rect 1626 438 1646 441
rect 442 428 566 431
rect 698 428 894 431
rect 906 428 1054 431
rect 1058 428 1222 431
rect 1490 428 1654 431
rect 1658 428 1918 431
rect 410 418 438 421
rect 514 418 630 421
rect 850 418 1654 421
rect 1658 418 1678 421
rect 1706 418 1710 421
rect 1746 418 1846 421
rect 1866 418 1870 421
rect 1906 418 1918 421
rect 650 408 750 411
rect 826 408 1190 411
rect 1554 408 1734 411
rect 496 403 498 407
rect 502 403 505 407
rect 510 403 512 407
rect 1528 403 1530 407
rect 1534 403 1537 407
rect 1542 403 1544 407
rect 578 398 622 401
rect 626 398 734 401
rect 738 398 830 401
rect 898 398 1062 401
rect 1098 398 1110 401
rect 1250 398 1398 401
rect 1626 398 1678 401
rect 122 388 134 391
rect 138 388 382 391
rect 690 388 846 391
rect 850 388 870 391
rect 874 388 1286 391
rect 1330 388 1542 391
rect 1610 388 1630 391
rect 1674 388 1958 391
rect 322 378 518 381
rect 618 378 1353 381
rect 1594 378 1622 381
rect 1698 378 1718 381
rect 1722 378 1817 381
rect 58 368 158 371
rect 202 368 286 371
rect 318 371 321 378
rect 1350 372 1353 378
rect 1814 372 1817 378
rect 318 368 358 371
rect 826 368 854 371
rect 858 368 982 371
rect 994 368 1006 371
rect 1090 368 1094 371
rect 1102 368 1118 371
rect 1138 368 1206 371
rect 1354 368 1366 371
rect 1650 368 1734 371
rect 1818 368 1838 371
rect 1842 368 1942 371
rect 374 362 377 368
rect 398 362 401 368
rect 750 362 753 368
rect 806 362 809 368
rect 162 358 166 361
rect 290 358 326 361
rect 330 358 374 361
rect 402 358 430 361
rect 466 358 478 361
rect 562 358 598 361
rect 602 358 638 361
rect 658 358 670 361
rect 1102 361 1105 368
rect 810 358 1105 361
rect 1362 358 1558 361
rect 1570 358 1742 361
rect 1746 358 1782 361
rect 1790 358 1894 361
rect 182 352 185 358
rect 646 352 649 358
rect 18 348 142 351
rect 146 348 174 351
rect 282 348 350 351
rect 402 348 406 351
rect 658 348 702 351
rect 714 348 774 351
rect 778 348 950 351
rect 986 348 1110 351
rect 1290 348 1302 351
rect 1306 348 1694 351
rect 1790 351 1793 358
rect 1778 348 1793 351
rect 1810 348 1889 351
rect 178 338 190 341
rect 194 338 294 341
rect 306 338 438 341
rect 490 338 494 341
rect 538 338 582 341
rect 618 338 662 341
rect 666 338 686 341
rect 722 338 838 341
rect 874 338 934 341
rect 974 341 977 348
rect 1886 342 1889 348
rect 974 338 998 341
rect 1058 338 1062 341
rect 1106 338 1134 341
rect 1138 338 1150 341
rect 1210 338 1278 341
rect 1338 338 1422 341
rect 1662 338 1694 341
rect 1662 332 1665 338
rect 106 328 158 331
rect 442 328 462 331
rect 466 328 574 331
rect 578 328 710 331
rect 762 328 798 331
rect 802 328 990 331
rect 994 328 1158 331
rect 1170 328 1430 331
rect 1790 331 1793 338
rect 1790 328 1846 331
rect 1978 328 2014 331
rect 74 318 126 321
rect 170 318 198 321
rect 298 318 334 321
rect 390 321 393 328
rect 390 318 470 321
rect 698 318 774 321
rect 786 318 806 321
rect 826 318 990 321
rect 1010 318 1038 321
rect 1050 318 1054 321
rect 1066 318 1126 321
rect 1306 318 1366 321
rect 1730 318 1766 321
rect 1770 318 1814 321
rect 290 308 542 311
rect 594 308 966 311
rect 1122 308 1422 311
rect 1426 308 1614 311
rect 1970 308 1974 311
rect 1016 303 1018 307
rect 1022 303 1025 307
rect 1030 303 1032 307
rect 418 298 502 301
rect 514 298 550 301
rect 554 298 614 301
rect 618 298 670 301
rect 674 298 718 301
rect 722 298 774 301
rect 778 298 830 301
rect 1154 298 1190 301
rect 1514 298 1574 301
rect 1802 298 1870 301
rect 314 288 342 291
rect 346 288 350 291
rect 466 288 822 291
rect 826 288 1078 291
rect 1082 288 1710 291
rect 1722 288 1790 291
rect 234 278 326 281
rect 442 278 494 281
rect 498 278 617 281
rect 634 278 814 281
rect 858 278 870 281
rect 882 278 934 281
rect 1218 278 1446 281
rect 1450 278 1598 281
rect 1634 278 1670 281
rect 1682 278 1878 281
rect 1882 278 1926 281
rect 358 271 361 278
rect 614 272 617 278
rect 258 268 361 271
rect 402 268 454 271
rect 458 268 478 271
rect 634 268 654 271
rect 658 268 694 271
rect 830 271 833 278
rect 950 272 953 278
rect 1046 272 1049 278
rect 1118 272 1121 278
rect 802 268 846 271
rect 866 268 902 271
rect 914 268 918 271
rect 930 268 942 271
rect 962 268 966 271
rect 1098 268 1118 271
rect 1138 268 1166 271
rect 1174 271 1177 278
rect 1174 268 1254 271
rect 1282 268 1334 271
rect 1406 268 1462 271
rect 1482 268 1558 271
rect 1562 268 1606 271
rect 1610 268 1798 271
rect 1818 268 1902 271
rect 1906 268 1982 271
rect 134 261 137 268
rect 558 262 561 268
rect 66 258 137 261
rect 226 258 326 261
rect 330 258 462 261
rect 546 258 550 261
rect 718 261 721 268
rect 766 262 769 268
rect 594 258 721 261
rect 730 258 734 261
rect 834 258 881 261
rect 890 258 894 261
rect 974 261 977 268
rect 938 258 977 261
rect 982 262 985 268
rect 1406 262 1409 268
rect 1002 258 1006 261
rect 1042 258 1134 261
rect 1146 258 1206 261
rect 1242 258 1246 261
rect 1274 258 1318 261
rect 1450 258 1566 261
rect 1642 258 1646 261
rect 1806 261 1809 268
rect 1762 258 1809 261
rect 1930 258 1998 261
rect 2002 258 2030 261
rect 878 252 881 258
rect 386 248 457 251
rect 490 248 502 251
rect 618 248 630 251
rect 654 248 705 251
rect 718 248 726 251
rect 730 248 742 251
rect 906 248 1126 251
rect 1130 248 1182 251
rect 1210 248 1222 251
rect 1226 248 1246 251
rect 1626 248 1638 251
rect 1682 248 1862 251
rect 1866 248 1942 251
rect 454 242 457 248
rect 654 242 657 248
rect 702 242 705 248
rect 778 238 1038 241
rect 1266 238 1302 241
rect 154 228 598 231
rect 610 228 622 231
rect 690 228 814 231
rect 1050 228 1062 231
rect 1194 228 1822 231
rect 626 218 662 221
rect 666 218 782 221
rect 874 218 897 221
rect 1182 221 1185 228
rect 946 218 1185 221
rect 1962 218 1990 221
rect 798 212 801 218
rect 894 212 897 218
rect 946 208 1006 211
rect 1162 208 1278 211
rect 1282 208 1294 211
rect 496 203 498 207
rect 502 203 505 207
rect 510 203 512 207
rect 1528 203 1530 207
rect 1534 203 1537 207
rect 1542 203 1544 207
rect 818 198 1142 201
rect 1994 198 1998 201
rect 374 188 382 191
rect 386 188 678 191
rect 698 188 886 191
rect 962 188 1638 191
rect 1954 188 1969 191
rect 1966 182 1969 188
rect 506 178 566 181
rect 1026 178 1422 181
rect 1426 178 1462 181
rect 1602 178 1606 181
rect 1610 178 1622 181
rect 1626 178 1782 181
rect 1786 178 1806 181
rect 318 172 321 178
rect 258 168 302 171
rect 346 168 518 171
rect 522 168 550 171
rect 658 168 678 171
rect 682 168 726 171
rect 890 168 1006 171
rect 1010 168 1110 171
rect 1154 168 1158 171
rect 1418 168 1462 171
rect 1466 168 1558 171
rect 1634 168 1686 171
rect 1690 168 1854 171
rect 1858 168 1870 171
rect 878 162 881 168
rect 106 158 118 161
rect 266 158 294 161
rect 298 158 862 161
rect 866 158 878 161
rect 1074 158 1150 161
rect 1178 158 1222 161
rect 1370 158 1654 161
rect 114 148 142 151
rect 146 148 182 151
rect 202 148 278 151
rect 322 148 342 151
rect 450 148 537 151
rect 618 148 793 151
rect 802 148 998 151
rect 1162 148 1190 151
rect 1362 148 1438 151
rect 1442 148 1550 151
rect 1554 148 1670 151
rect 1674 148 1694 151
rect 1738 148 1830 151
rect 1834 148 1862 151
rect 534 142 537 148
rect 98 138 150 141
rect 266 138 318 141
rect 322 138 326 141
rect 370 138 382 141
rect 386 138 430 141
rect 722 138 726 141
rect 790 141 793 148
rect 790 138 822 141
rect 1186 138 1190 141
rect 1434 138 1462 141
rect 1466 138 1598 141
rect 1658 138 1678 141
rect 58 128 110 131
rect 362 128 390 131
rect 402 128 414 131
rect 746 128 790 131
rect 982 131 985 138
rect 982 128 990 131
rect 1106 128 1142 131
rect 1254 131 1257 138
rect 1630 132 1633 138
rect 1146 128 1257 131
rect 1446 128 1510 131
rect 1446 122 1449 128
rect 394 118 574 121
rect 1106 118 1206 121
rect 1866 118 1870 121
rect 262 112 265 118
rect 266 108 286 111
rect 690 108 846 111
rect 1642 108 1734 111
rect 1738 108 1766 111
rect 1016 103 1018 107
rect 1022 103 1025 107
rect 1030 103 1032 107
rect 250 98 758 101
rect 842 98 862 101
rect 866 98 910 101
rect 1578 98 1622 101
rect 1994 98 2014 101
rect 290 88 414 91
rect 418 88 878 91
rect 1034 88 1038 91
rect 1042 88 1118 91
rect 1154 88 1190 91
rect 1194 88 1222 91
rect 1314 88 1334 91
rect 1338 88 1374 91
rect 1538 88 1566 91
rect 1594 88 1614 91
rect 1986 88 2022 91
rect 298 78 686 81
rect 786 78 806 81
rect 1082 78 1166 81
rect 18 68 30 71
rect 34 68 70 71
rect 142 68 313 71
rect 702 71 705 78
rect 1214 72 1217 78
rect 602 68 846 71
rect 850 68 918 71
rect 922 68 942 71
rect 946 68 1054 71
rect 1178 68 1214 71
rect 1310 71 1313 78
rect 1310 68 1374 71
rect 1606 71 1609 78
rect 1718 71 1721 78
rect 1606 68 1766 71
rect 1770 68 1862 71
rect 142 62 145 68
rect 158 62 161 68
rect 310 62 313 68
rect 194 58 270 61
rect 290 58 294 61
rect 314 58 438 61
rect 442 58 470 61
rect 586 58 654 61
rect 866 58 958 61
rect 1086 61 1089 68
rect 1086 58 1134 61
rect 1170 58 1214 61
rect 2026 58 2046 61
rect 2078 61 2082 62
rect 2050 58 2082 61
rect 414 48 486 51
rect 666 48 678 51
rect 682 48 782 51
rect 786 48 1126 51
rect 1130 48 1158 51
rect 1210 48 1270 51
rect 414 42 417 48
rect 1994 8 1998 11
rect 2018 8 2030 11
rect 496 3 498 7
rect 502 3 505 7
rect 510 3 512 7
rect 1528 3 1530 7
rect 1534 3 1537 7
rect 1542 3 1544 7
<< m4contact >>
rect -26 1818 -22 1822
rect 498 1803 502 1807
rect 506 1803 509 1807
rect 509 1803 510 1807
rect 1530 1803 1534 1807
rect 1538 1803 1541 1807
rect 1541 1803 1542 1807
rect 6 1798 10 1802
rect 22 1788 26 1792
rect 6 1778 10 1782
rect 1966 1768 1970 1772
rect 1934 1758 1938 1762
rect 1670 1738 1674 1742
rect 1966 1728 1970 1732
rect 1118 1718 1122 1722
rect 1902 1718 1906 1722
rect 1018 1703 1022 1707
rect 1026 1703 1029 1707
rect 1029 1703 1030 1707
rect 486 1698 490 1702
rect 1062 1678 1066 1682
rect 1550 1668 1554 1672
rect 1902 1668 1906 1672
rect 1126 1658 1130 1662
rect 2014 1658 2018 1662
rect 662 1648 666 1652
rect 718 1638 722 1642
rect 1974 1638 1978 1642
rect 734 1628 738 1632
rect 246 1618 250 1622
rect 1230 1618 1234 1622
rect 498 1603 502 1607
rect 506 1603 509 1607
rect 509 1603 510 1607
rect 1530 1603 1534 1607
rect 1538 1603 1541 1607
rect 1541 1603 1542 1607
rect 774 1598 778 1602
rect 1694 1598 1698 1602
rect 30 1588 34 1592
rect 846 1588 850 1592
rect 630 1578 634 1582
rect 214 1558 218 1562
rect 1934 1558 1938 1562
rect 1062 1548 1066 1552
rect 1118 1548 1122 1552
rect 446 1538 450 1542
rect 1518 1538 1522 1542
rect 1902 1538 1906 1542
rect 142 1528 146 1532
rect 1382 1528 1386 1532
rect 1750 1528 1754 1532
rect 614 1508 618 1512
rect 1966 1508 1970 1512
rect 1018 1503 1022 1507
rect 1026 1503 1029 1507
rect 1029 1503 1030 1507
rect 390 1498 394 1502
rect 750 1498 754 1502
rect 1254 1498 1258 1502
rect 1822 1498 1826 1502
rect 1838 1498 1842 1502
rect 622 1488 626 1492
rect 1694 1488 1698 1492
rect 254 1478 258 1482
rect 630 1478 634 1482
rect 846 1478 850 1482
rect 1238 1468 1242 1472
rect 1742 1468 1746 1472
rect 246 1458 250 1462
rect 542 1458 546 1462
rect 1550 1458 1554 1462
rect 1854 1458 1858 1462
rect 126 1448 130 1452
rect 1054 1448 1058 1452
rect 1206 1448 1210 1452
rect 1710 1448 1714 1452
rect 1830 1448 1834 1452
rect 1902 1448 1906 1452
rect 134 1438 138 1442
rect 190 1438 194 1442
rect 2014 1448 2018 1452
rect 1854 1438 1858 1442
rect 222 1428 226 1432
rect 1006 1428 1010 1432
rect 1230 1428 1234 1432
rect 1278 1428 1282 1432
rect 1998 1428 2002 1432
rect 678 1418 682 1422
rect 1158 1418 1162 1422
rect 1614 1418 1618 1422
rect 1958 1418 1962 1422
rect 926 1408 930 1412
rect 1286 1408 1290 1412
rect 1470 1408 1474 1412
rect 1734 1408 1738 1412
rect 1998 1408 2002 1412
rect 498 1403 502 1407
rect 506 1403 509 1407
rect 509 1403 510 1407
rect 1530 1403 1534 1407
rect 1538 1403 1541 1407
rect 1541 1403 1542 1407
rect 1734 1398 1738 1402
rect 214 1388 218 1392
rect 1078 1388 1082 1392
rect 1278 1388 1282 1392
rect 2022 1378 2026 1382
rect 1270 1368 1274 1372
rect 1646 1368 1650 1372
rect 2030 1368 2034 1372
rect 134 1358 138 1362
rect 918 1358 922 1362
rect 958 1358 962 1362
rect 1206 1358 1210 1362
rect 1254 1358 1258 1362
rect 1990 1358 1994 1362
rect 190 1348 194 1352
rect 662 1348 666 1352
rect 1230 1348 1234 1352
rect 1374 1348 1378 1352
rect 390 1338 394 1342
rect 526 1338 530 1342
rect 1286 1338 1290 1342
rect 1518 1338 1522 1342
rect 1790 1338 1794 1342
rect 1974 1338 1978 1342
rect 806 1328 810 1332
rect 1654 1328 1658 1332
rect 398 1318 402 1322
rect 670 1318 674 1322
rect 822 1318 826 1322
rect 998 1318 1002 1322
rect 1358 1318 1362 1322
rect 414 1308 418 1312
rect 438 1308 442 1312
rect 758 1308 762 1312
rect 1150 1308 1154 1312
rect 1018 1303 1022 1307
rect 1026 1303 1029 1307
rect 1029 1303 1030 1307
rect 1966 1298 1970 1302
rect 1982 1298 1986 1302
rect 486 1288 490 1292
rect 502 1288 506 1292
rect 894 1288 898 1292
rect 1094 1288 1098 1292
rect 1558 1288 1562 1292
rect 1758 1288 1762 1292
rect 1822 1288 1826 1292
rect 1894 1288 1898 1292
rect 2046 1288 2050 1292
rect 406 1278 410 1282
rect 830 1278 834 1282
rect 846 1278 850 1282
rect 870 1278 874 1282
rect 1158 1278 1162 1282
rect 2022 1278 2026 1282
rect 470 1268 474 1272
rect 582 1268 586 1272
rect 662 1268 666 1272
rect 1038 1268 1042 1272
rect 1062 1268 1066 1272
rect 1390 1268 1394 1272
rect 1590 1268 1594 1272
rect 1686 1268 1690 1272
rect 2046 1268 2050 1272
rect 126 1258 130 1262
rect 342 1258 346 1262
rect 1398 1258 1402 1262
rect 1614 1258 1618 1262
rect 1742 1258 1746 1262
rect 1838 1248 1842 1252
rect 374 1238 378 1242
rect 438 1238 442 1242
rect 1134 1238 1138 1242
rect 1710 1238 1714 1242
rect 1718 1238 1722 1242
rect 1726 1238 1730 1242
rect 534 1228 538 1232
rect 766 1218 770 1222
rect 1630 1218 1634 1222
rect 1886 1218 1890 1222
rect 1910 1218 1914 1222
rect 814 1208 818 1212
rect 1734 1208 1738 1212
rect 498 1203 502 1207
rect 506 1203 509 1207
rect 509 1203 510 1207
rect 1530 1203 1534 1207
rect 1538 1203 1541 1207
rect 1541 1203 1542 1207
rect 1598 1198 1602 1202
rect 646 1178 650 1182
rect 862 1178 866 1182
rect 582 1168 586 1172
rect 654 1158 658 1162
rect 926 1158 930 1162
rect 1190 1158 1194 1162
rect 1454 1158 1458 1162
rect 1574 1158 1578 1162
rect 422 1148 426 1152
rect 998 1148 1002 1152
rect 1054 1148 1058 1152
rect 1294 1148 1298 1152
rect 1382 1148 1386 1152
rect 1510 1148 1514 1152
rect 1606 1148 1610 1152
rect 542 1138 546 1142
rect 1174 1138 1178 1142
rect 1310 1138 1314 1142
rect 1646 1138 1650 1142
rect 678 1128 682 1132
rect 1158 1128 1162 1132
rect 1462 1128 1466 1132
rect 1638 1128 1642 1132
rect 1750 1128 1754 1132
rect 1942 1118 1946 1122
rect 486 1108 490 1112
rect 1286 1108 1290 1112
rect 1018 1103 1022 1107
rect 1026 1103 1029 1107
rect 1029 1103 1030 1107
rect 710 1098 714 1102
rect 726 1098 730 1102
rect 1510 1098 1514 1102
rect 1934 1098 1938 1102
rect 414 1088 418 1092
rect 1726 1088 1730 1092
rect 254 1078 258 1082
rect 310 1078 314 1082
rect 398 1078 402 1082
rect 414 1078 418 1082
rect 646 1078 650 1082
rect 686 1078 690 1082
rect 726 1078 730 1082
rect 1294 1078 1298 1082
rect 1662 1078 1666 1082
rect 1702 1078 1706 1082
rect 174 1068 178 1072
rect 542 1068 546 1072
rect 574 1068 578 1072
rect 670 1068 674 1072
rect 926 1068 930 1072
rect 1470 1068 1474 1072
rect 1654 1068 1658 1072
rect 414 1058 418 1062
rect 422 1058 426 1062
rect 430 1058 434 1062
rect 686 1058 690 1062
rect 958 1058 962 1062
rect 1238 1058 1242 1062
rect 1718 1058 1722 1062
rect 1926 1058 1930 1062
rect 318 1048 322 1052
rect 694 1048 698 1052
rect 854 1048 858 1052
rect 1798 1048 1802 1052
rect 2038 1048 2042 1052
rect 214 1038 218 1042
rect 438 1038 442 1042
rect 1126 1038 1130 1042
rect 1214 1038 1218 1042
rect 1134 1028 1138 1032
rect 1166 1028 1170 1032
rect 2006 1028 2010 1032
rect 806 1018 810 1022
rect 1486 1018 1490 1022
rect 894 1008 898 1012
rect 1910 1008 1914 1012
rect 498 1003 502 1007
rect 506 1003 509 1007
rect 509 1003 510 1007
rect 1530 1003 1534 1007
rect 1538 1003 1541 1007
rect 1541 1003 1542 1007
rect 766 998 770 1002
rect 30 988 34 992
rect 406 988 410 992
rect 622 988 626 992
rect 870 988 874 992
rect 1694 988 1698 992
rect 758 978 762 982
rect 862 978 866 982
rect 926 978 930 982
rect 534 968 538 972
rect 726 968 730 972
rect 742 968 746 972
rect 1262 968 1266 972
rect 1622 968 1626 972
rect 222 958 226 962
rect 398 958 402 962
rect 470 958 474 962
rect 646 948 650 952
rect 734 948 738 952
rect 830 948 834 952
rect 1390 948 1394 952
rect 1454 948 1458 952
rect 1462 948 1466 952
rect 462 938 466 942
rect 478 938 482 942
rect 598 938 602 942
rect 638 938 642 942
rect 798 938 802 942
rect 822 938 826 942
rect 998 938 1002 942
rect 1502 938 1506 942
rect 1622 938 1626 942
rect 1654 938 1658 942
rect 406 928 410 932
rect 854 928 858 932
rect 902 928 906 932
rect 1542 928 1546 932
rect 1590 928 1594 932
rect 310 918 314 922
rect 806 918 810 922
rect 1158 918 1162 922
rect 374 908 378 912
rect 758 908 762 912
rect 1046 908 1050 912
rect 1598 908 1602 912
rect 1018 903 1022 907
rect 1026 903 1029 907
rect 1029 903 1030 907
rect 326 888 330 892
rect 606 888 610 892
rect 654 888 658 892
rect 702 888 706 892
rect 838 888 842 892
rect 846 888 850 892
rect 1046 888 1050 892
rect 1150 888 1154 892
rect 1478 888 1482 892
rect 1598 888 1602 892
rect 654 878 658 882
rect 446 868 450 872
rect 990 868 994 872
rect 1062 868 1066 872
rect 1702 868 1706 872
rect 1766 868 1770 872
rect 126 858 130 862
rect 134 858 138 862
rect 750 858 754 862
rect 782 858 786 862
rect 822 858 826 862
rect 870 858 874 862
rect 1438 858 1442 862
rect 1910 858 1914 862
rect 1950 858 1954 862
rect 2014 858 2018 862
rect 686 848 690 852
rect 790 848 794 852
rect 1006 848 1010 852
rect 1622 848 1626 852
rect 1662 848 1666 852
rect 606 838 610 842
rect 1590 838 1594 842
rect 582 828 586 832
rect 622 828 626 832
rect 1686 828 1690 832
rect 614 818 618 822
rect 950 818 954 822
rect 1630 818 1634 822
rect 134 808 138 812
rect 182 808 186 812
rect 470 808 474 812
rect 830 808 834 812
rect 498 803 502 807
rect 506 803 509 807
rect 509 803 510 807
rect 1530 803 1534 807
rect 1538 803 1541 807
rect 1541 803 1542 807
rect 958 798 962 802
rect 774 788 778 792
rect 1158 788 1162 792
rect 1190 788 1194 792
rect 694 778 698 782
rect 1006 778 1010 782
rect 1190 778 1194 782
rect 526 768 530 772
rect 726 768 730 772
rect 990 768 994 772
rect 1406 768 1410 772
rect 1606 768 1610 772
rect 470 758 474 762
rect 494 758 498 762
rect 710 758 714 762
rect 750 758 754 762
rect 1070 758 1074 762
rect 1150 758 1154 762
rect 1582 758 1586 762
rect 1614 758 1618 762
rect 550 748 554 752
rect 590 748 594 752
rect 142 738 146 742
rect 182 738 186 742
rect 726 748 730 752
rect 742 748 746 752
rect 766 748 770 752
rect 846 748 850 752
rect 886 748 890 752
rect 1054 748 1058 752
rect 1062 748 1066 752
rect 1294 748 1298 752
rect 1598 748 1602 752
rect 1942 748 1946 752
rect 670 738 674 742
rect 734 738 738 742
rect 750 738 754 742
rect 774 738 778 742
rect 830 738 834 742
rect 918 738 922 742
rect 1238 738 1242 742
rect 1438 738 1442 742
rect 1542 738 1546 742
rect 1702 738 1706 742
rect 174 728 178 732
rect 718 728 722 732
rect 782 728 786 732
rect 846 728 850 732
rect 1110 728 1114 732
rect 1294 728 1298 732
rect 1422 728 1426 732
rect 1446 728 1450 732
rect 1638 728 1642 732
rect 1694 728 1698 732
rect 1934 728 1938 732
rect 326 718 330 722
rect 694 718 698 722
rect 1166 718 1170 722
rect 1222 718 1226 722
rect 1806 718 1810 722
rect 286 708 290 712
rect 1018 703 1022 707
rect 1026 703 1029 707
rect 1029 703 1030 707
rect 566 698 570 702
rect 758 698 762 702
rect 1510 698 1514 702
rect 574 688 578 692
rect 982 688 986 692
rect 462 678 466 682
rect 1190 678 1194 682
rect 1350 678 1354 682
rect 1470 678 1474 682
rect 1678 678 1682 682
rect 2014 678 2018 682
rect 486 668 490 672
rect 518 668 522 672
rect 638 668 642 672
rect 854 668 858 672
rect 926 668 930 672
rect 998 668 1002 672
rect 1286 668 1290 672
rect 1494 668 1498 672
rect 1526 668 1530 672
rect 1662 668 1666 672
rect 142 658 146 662
rect 286 658 290 662
rect 566 658 570 662
rect 702 658 706 662
rect 814 658 818 662
rect 1614 658 1618 662
rect 1646 658 1650 662
rect 1686 658 1690 662
rect 1934 658 1938 662
rect 1950 658 1954 662
rect 2014 658 2018 662
rect 550 648 554 652
rect 958 648 962 652
rect 1270 648 1274 652
rect 886 638 890 642
rect 934 638 938 642
rect 1238 628 1242 632
rect 838 618 842 622
rect 902 618 906 622
rect 1262 618 1266 622
rect 1358 618 1362 622
rect 1390 608 1394 612
rect 498 603 502 607
rect 506 603 509 607
rect 509 603 510 607
rect 1530 603 1534 607
rect 1538 603 1541 607
rect 1541 603 1542 607
rect 262 588 266 592
rect 686 588 690 592
rect 1038 588 1042 592
rect 1182 588 1186 592
rect 1486 588 1490 592
rect 790 578 794 582
rect 350 568 354 572
rect 1102 568 1106 572
rect 1166 568 1170 572
rect 2006 568 2010 572
rect 342 558 346 562
rect 406 558 410 562
rect 582 558 586 562
rect 878 558 882 562
rect 1646 558 1650 562
rect 590 548 594 552
rect 1190 548 1194 552
rect 1886 548 1890 552
rect 598 538 602 542
rect 630 538 634 542
rect 1118 538 1122 542
rect 1174 538 1178 542
rect 1934 538 1938 542
rect 678 528 682 532
rect 702 528 706 532
rect 998 528 1002 532
rect 1638 528 1642 532
rect 2022 528 2026 532
rect 1046 518 1050 522
rect 1174 518 1178 522
rect 2038 518 2042 522
rect 126 508 130 512
rect 598 508 602 512
rect 1086 508 1090 512
rect 1142 508 1146 512
rect 2046 508 2050 512
rect 1018 503 1022 507
rect 1026 503 1029 507
rect 1029 503 1030 507
rect 726 498 730 502
rect 902 498 906 502
rect 1046 498 1050 502
rect 1926 498 1930 502
rect 870 488 874 492
rect 918 488 922 492
rect 2038 488 2042 492
rect 222 478 226 482
rect 318 478 322 482
rect 1486 478 1490 482
rect 2014 478 2018 482
rect 30 468 34 472
rect 494 468 498 472
rect 1038 468 1042 472
rect 1054 468 1058 472
rect 1062 468 1066 472
rect 1086 468 1090 472
rect 1134 468 1138 472
rect 1478 468 1482 472
rect 1550 468 1554 472
rect 2022 468 2026 472
rect 2038 468 2042 472
rect 126 458 130 462
rect 862 458 866 462
rect 966 458 970 462
rect 982 458 986 462
rect 1006 458 1010 462
rect 1166 458 1170 462
rect 1494 458 1498 462
rect 1958 458 1962 462
rect 494 448 498 452
rect 894 448 898 452
rect 998 448 1002 452
rect 1158 448 1162 452
rect 1270 448 1274 452
rect 1278 448 1282 452
rect 1494 448 1498 452
rect 1646 448 1650 452
rect 518 438 522 442
rect 1086 438 1090 442
rect 1622 438 1626 442
rect 902 428 906 432
rect 438 418 442 422
rect 630 418 634 422
rect 846 418 850 422
rect 1654 418 1658 422
rect 1710 418 1714 422
rect 1870 418 1874 422
rect 1902 418 1906 422
rect 646 408 650 412
rect 1190 408 1194 412
rect 1550 408 1554 412
rect 498 403 502 407
rect 506 403 509 407
rect 509 403 510 407
rect 1530 403 1534 407
rect 1538 403 1541 407
rect 1541 403 1542 407
rect 622 398 626 402
rect 1062 398 1066 402
rect 1094 398 1098 402
rect 286 368 290 372
rect 398 368 402 372
rect 750 368 754 372
rect 822 368 826 372
rect 982 368 986 372
rect 1086 368 1090 372
rect 1134 368 1138 372
rect 1646 368 1650 372
rect 166 358 170 362
rect 374 358 378 362
rect 806 358 810 362
rect 1566 358 1570 362
rect 174 348 178 352
rect 182 348 186 352
rect 398 348 402 352
rect 646 348 650 352
rect 702 348 706 352
rect 710 348 714 352
rect 950 348 954 352
rect 982 348 986 352
rect 294 338 298 342
rect 494 338 498 342
rect 614 338 618 342
rect 718 338 722 342
rect 1062 338 1066 342
rect 1206 338 1210 342
rect 438 328 442 332
rect 710 328 714 332
rect 1166 328 1170 332
rect 1974 328 1978 332
rect 294 318 298 322
rect 774 318 778 322
rect 1046 318 1050 322
rect 966 308 970 312
rect 1966 308 1970 312
rect 1018 303 1022 307
rect 1026 303 1029 307
rect 1029 303 1030 307
rect 502 298 506 302
rect 1150 298 1154 302
rect 1798 298 1802 302
rect 350 288 354 292
rect 1710 288 1714 292
rect 1718 288 1722 292
rect 814 278 818 282
rect 934 278 938 282
rect 1046 278 1050 282
rect 1174 278 1178 282
rect 630 268 634 272
rect 902 268 906 272
rect 918 268 922 272
rect 926 268 930 272
rect 950 268 954 272
rect 958 268 962 272
rect 1118 268 1122 272
rect 1798 268 1802 272
rect 542 258 546 262
rect 558 258 562 262
rect 726 258 730 262
rect 766 258 770 262
rect 982 258 986 262
rect 998 258 1002 262
rect 1038 258 1042 262
rect 1142 258 1146 262
rect 1238 258 1242 262
rect 1638 258 1642 262
rect 1998 258 2002 262
rect 614 248 618 252
rect 1182 248 1186 252
rect 1222 248 1226 252
rect 1862 248 1866 252
rect 1038 238 1042 242
rect 1262 238 1266 242
rect 798 218 802 222
rect 1278 208 1282 212
rect 498 203 502 207
rect 506 203 509 207
rect 509 203 510 207
rect 1530 203 1534 207
rect 1538 203 1541 207
rect 1541 203 1542 207
rect 1142 198 1146 202
rect 1990 198 1994 202
rect 886 188 890 192
rect 318 178 322 182
rect 1606 178 1610 182
rect 654 168 658 172
rect 878 168 882 172
rect 886 168 890 172
rect 1110 168 1114 172
rect 1158 168 1162 172
rect 1070 158 1074 162
rect 182 148 186 152
rect 1670 148 1674 152
rect 718 138 722 142
rect 1190 138 1194 142
rect 1630 138 1634 142
rect 1102 128 1106 132
rect 262 118 266 122
rect 846 108 850 112
rect 1638 108 1642 112
rect 1018 103 1022 107
rect 1026 103 1029 107
rect 1029 103 1030 107
rect 862 98 866 102
rect 1574 98 1578 102
rect 286 88 290 92
rect 1150 88 1154 92
rect 294 78 298 82
rect 30 68 34 72
rect 1214 68 1218 72
rect 294 58 298 62
rect 2046 58 2050 62
rect 1998 8 2002 12
rect 2030 8 2034 12
rect 498 3 502 7
rect 506 3 509 7
rect 509 3 510 7
rect 1530 3 1534 7
rect 1538 3 1541 7
rect 1541 3 1542 7
<< metal4 >>
rect -22 1818 -18 1821
rect 496 1803 498 1807
rect 502 1803 505 1807
rect 510 1803 512 1807
rect 1528 1803 1530 1807
rect 1534 1803 1537 1807
rect 1542 1803 1544 1807
rect 6 1782 9 1798
rect 22 1792 25 1798
rect 1016 1703 1018 1707
rect 1022 1703 1025 1707
rect 1030 1703 1032 1707
rect 30 992 33 1588
rect 126 1262 129 1448
rect 134 1362 137 1438
rect 30 472 33 988
rect 134 862 137 1358
rect 126 512 129 858
rect 134 661 137 808
rect 142 742 145 1528
rect 190 1352 193 1438
rect 214 1392 217 1558
rect 246 1462 249 1618
rect 182 1348 190 1351
rect 174 732 177 1068
rect 182 812 185 1348
rect 182 672 185 738
rect 134 658 142 661
rect 30 72 33 468
rect 126 462 129 508
rect 158 361 161 368
rect 158 358 166 361
rect 182 352 185 668
rect 214 372 217 1038
rect 222 962 225 1428
rect 254 1082 257 1478
rect 390 1342 393 1498
rect 222 482 225 958
rect 310 922 313 1078
rect 318 1052 321 1058
rect 326 722 329 888
rect 286 662 289 708
rect 174 262 177 348
rect 182 152 185 348
rect 262 122 265 588
rect 342 571 345 1258
rect 374 912 377 1238
rect 398 1082 401 1318
rect 398 962 401 1078
rect 406 992 409 1278
rect 414 1092 417 1308
rect 438 1292 441 1308
rect 414 1062 417 1078
rect 422 1062 425 1148
rect 430 1062 433 1068
rect 438 1042 441 1238
rect 342 568 350 571
rect 286 92 289 368
rect 294 342 297 348
rect 294 82 297 318
rect 318 182 321 478
rect 342 291 345 558
rect 398 372 401 958
rect 406 562 409 928
rect 446 872 449 1538
rect 486 1292 489 1698
rect 496 1603 498 1607
rect 502 1603 505 1607
rect 510 1603 512 1607
rect 496 1403 498 1407
rect 502 1403 505 1407
rect 510 1403 512 1407
rect 498 1288 502 1291
rect 470 1262 473 1268
rect 496 1203 498 1207
rect 502 1203 505 1207
rect 510 1203 512 1207
rect 462 682 465 938
rect 470 812 473 958
rect 478 942 481 948
rect 470 762 473 808
rect 486 672 489 1108
rect 496 1003 498 1007
rect 502 1003 505 1007
rect 510 1003 512 1007
rect 496 803 498 807
rect 502 803 505 807
rect 510 803 512 807
rect 526 772 529 1338
rect 534 972 537 1228
rect 542 1142 545 1458
rect 586 1268 590 1271
rect 498 758 502 761
rect 496 603 498 607
rect 502 603 505 607
rect 510 603 512 607
rect 494 452 497 468
rect 518 442 521 668
rect 378 358 382 361
rect 402 348 406 351
rect 438 332 441 418
rect 496 403 498 407
rect 502 403 505 407
rect 510 403 512 407
rect 490 338 494 341
rect 342 288 350 291
rect 502 252 505 298
rect 542 262 545 1068
rect 550 652 553 748
rect 566 702 569 728
rect 574 692 577 1068
rect 582 832 585 1168
rect 594 938 598 941
rect 606 842 609 888
rect 566 442 569 658
rect 582 562 585 828
rect 614 822 617 1508
rect 622 992 625 1488
rect 630 1482 633 1578
rect 662 1352 665 1648
rect 662 1272 665 1288
rect 646 1082 649 1178
rect 638 932 641 938
rect 590 552 593 748
rect 598 512 601 538
rect 622 402 625 828
rect 634 668 638 671
rect 634 538 638 541
rect 614 342 617 358
rect 630 272 633 418
rect 646 412 649 948
rect 654 892 657 1158
rect 670 1072 673 1318
rect 678 1132 681 1418
rect 718 1101 721 1638
rect 714 1098 721 1101
rect 726 1082 729 1098
rect 690 1078 697 1081
rect 686 1012 689 1058
rect 694 1052 697 1078
rect 646 352 649 408
rect 554 258 558 261
rect 610 248 614 251
rect 496 203 498 207
rect 502 203 505 207
rect 510 203 512 207
rect 654 172 657 878
rect 674 738 681 741
rect 678 532 681 738
rect 686 592 689 848
rect 694 722 697 778
rect 702 662 705 888
rect 726 772 729 968
rect 734 952 737 1628
rect 714 758 718 761
rect 742 752 745 968
rect 750 862 753 1498
rect 762 1308 769 1311
rect 766 1222 769 1308
rect 758 952 761 978
rect 750 752 753 758
rect 718 732 721 748
rect 702 532 705 658
rect 702 352 705 528
rect 726 502 729 748
rect 738 738 742 741
rect 750 372 753 738
rect 758 702 761 908
rect 766 752 769 998
rect 774 792 777 1598
rect 846 1482 849 1588
rect 1062 1552 1065 1678
rect 1118 1552 1121 1718
rect 1016 1503 1018 1507
rect 1022 1503 1025 1507
rect 1030 1503 1032 1507
rect 806 1022 809 1328
rect 818 1318 822 1321
rect 894 1282 897 1288
rect 834 1278 838 1281
rect 866 1278 870 1281
rect 782 852 785 858
rect 778 738 782 741
rect 778 728 782 731
rect 702 302 705 348
rect 710 332 713 348
rect 718 142 721 338
rect 774 322 777 718
rect 790 582 793 848
rect 726 262 729 268
rect 770 258 774 261
rect 798 222 801 938
rect 806 362 809 918
rect 814 662 817 1208
rect 822 862 825 938
rect 830 812 833 948
rect 846 892 849 1278
rect 854 932 857 1048
rect 862 982 865 1178
rect 826 738 830 741
rect 838 622 841 888
rect 870 862 873 988
rect 846 732 849 748
rect 850 668 854 671
rect 870 522 873 858
rect 882 748 886 751
rect 870 492 873 518
rect 818 368 822 371
rect 818 278 822 281
rect 846 112 849 418
rect 862 102 865 458
rect 878 172 881 558
rect 886 462 889 638
rect 894 452 897 1008
rect 918 981 921 1358
rect 926 1162 929 1408
rect 930 1068 934 1071
rect 958 1062 961 1358
rect 994 1318 998 1321
rect 918 978 926 981
rect 998 942 1001 1148
rect 902 722 905 928
rect 910 738 918 741
rect 910 732 913 738
rect 926 662 929 668
rect 934 642 937 938
rect 994 868 998 871
rect 1006 852 1009 1428
rect 1016 1303 1018 1307
rect 1022 1303 1025 1307
rect 1030 1303 1032 1307
rect 1016 1103 1018 1107
rect 1022 1103 1025 1107
rect 1030 1103 1032 1107
rect 1016 903 1018 907
rect 1022 903 1025 907
rect 1030 903 1032 907
rect 902 502 905 618
rect 914 488 918 491
rect 902 272 905 428
rect 950 352 953 818
rect 958 652 961 798
rect 990 691 993 768
rect 986 688 993 691
rect 998 672 1001 688
rect 938 278 942 281
rect 918 272 921 278
rect 950 272 953 348
rect 958 342 961 648
rect 974 461 977 468
rect 974 458 982 461
rect 958 272 961 338
rect 966 312 969 458
rect 998 452 1001 528
rect 1006 462 1009 778
rect 1016 703 1018 707
rect 1022 703 1025 707
rect 1030 703 1032 707
rect 1038 592 1041 1268
rect 1054 1152 1057 1448
rect 1062 1262 1065 1268
rect 1046 912 1049 1008
rect 1046 522 1049 888
rect 1058 868 1062 871
rect 1016 503 1018 507
rect 1022 503 1025 507
rect 1030 503 1032 507
rect 1046 472 1049 498
rect 1054 472 1057 748
rect 1062 742 1065 748
rect 982 352 985 368
rect 926 262 929 268
rect 982 262 985 348
rect 1016 303 1018 307
rect 1022 303 1025 307
rect 1030 303 1032 307
rect 1006 261 1009 298
rect 1002 258 1009 261
rect 1038 262 1041 468
rect 1046 322 1049 458
rect 1062 402 1065 468
rect 1058 338 1062 341
rect 1046 282 1049 288
rect 1038 242 1041 258
rect 886 172 889 188
rect 1070 162 1073 758
rect 1078 502 1081 1388
rect 1094 1282 1097 1288
rect 1126 1042 1129 1658
rect 1134 1032 1137 1238
rect 1150 892 1153 1308
rect 1158 1282 1161 1418
rect 1206 1362 1209 1448
rect 1230 1432 1233 1618
rect 1528 1603 1530 1607
rect 1534 1603 1537 1607
rect 1542 1603 1544 1607
rect 1226 1348 1230 1351
rect 1158 1132 1161 1278
rect 1178 1138 1182 1141
rect 1158 922 1161 1128
rect 1150 762 1153 888
rect 1086 482 1089 508
rect 1086 442 1089 468
rect 1094 402 1097 498
rect 1090 368 1094 371
rect 1102 132 1105 568
rect 1110 172 1113 728
rect 1118 272 1121 538
rect 1150 511 1153 518
rect 1146 508 1153 511
rect 1134 472 1137 488
rect 1130 368 1134 371
rect 1150 302 1153 508
rect 1158 452 1161 788
rect 1166 722 1169 1028
rect 1190 792 1193 1158
rect 1238 1062 1241 1468
rect 1254 1362 1257 1498
rect 1278 1392 1281 1428
rect 1190 682 1193 778
rect 1166 462 1169 568
rect 1174 522 1177 538
rect 1166 332 1169 338
rect 1174 272 1177 278
rect 1142 202 1145 258
rect 1182 252 1185 588
rect 1190 412 1193 548
rect 1150 168 1158 171
rect 1016 103 1018 107
rect 1022 103 1025 107
rect 1030 103 1032 107
rect 1150 92 1153 168
rect 1190 142 1193 408
rect 1206 342 1209 538
rect 294 62 297 78
rect 1214 72 1217 1038
rect 1222 252 1225 718
rect 1238 632 1241 738
rect 1262 622 1265 968
rect 1270 652 1273 1368
rect 1286 1342 1289 1408
rect 1370 1348 1374 1351
rect 1286 1112 1289 1338
rect 1358 1302 1361 1318
rect 1382 1152 1385 1528
rect 1294 1082 1297 1148
rect 1306 1138 1310 1141
rect 1390 952 1393 1268
rect 1390 872 1393 948
rect 1294 732 1297 748
rect 1346 678 1350 681
rect 1286 672 1289 678
rect 1358 622 1361 658
rect 1390 612 1393 868
rect 1398 771 1401 1258
rect 1454 952 1457 1158
rect 1462 952 1465 1128
rect 1470 1072 1473 1408
rect 1518 1342 1521 1538
rect 1550 1462 1553 1668
rect 1528 1403 1530 1407
rect 1534 1403 1537 1407
rect 1542 1403 1544 1407
rect 1510 1102 1513 1148
rect 1442 858 1446 861
rect 1398 768 1406 771
rect 1442 738 1446 741
rect 1422 732 1425 738
rect 1442 728 1446 731
rect 1466 678 1470 681
rect 1478 472 1481 888
rect 1486 592 1489 1018
rect 1506 938 1513 941
rect 1510 702 1513 938
rect 1518 671 1521 1298
rect 1554 1288 1558 1291
rect 1586 1268 1590 1271
rect 1614 1262 1617 1418
rect 1528 1203 1530 1207
rect 1534 1203 1537 1207
rect 1542 1203 1544 1207
rect 1528 1003 1530 1007
rect 1534 1003 1537 1007
rect 1542 1003 1544 1007
rect 1538 928 1542 931
rect 1528 803 1530 807
rect 1534 803 1537 807
rect 1542 803 1544 807
rect 1546 738 1550 741
rect 1518 668 1526 671
rect 1486 482 1489 488
rect 1494 462 1497 668
rect 1528 603 1530 607
rect 1534 603 1537 607
rect 1542 603 1544 607
rect 1494 452 1497 458
rect 1262 448 1270 451
rect 1242 258 1246 261
rect 1262 242 1265 448
rect 1278 212 1281 448
rect 1550 412 1553 468
rect 1528 403 1530 407
rect 1534 403 1537 407
rect 1542 403 1544 407
rect 1566 362 1569 438
rect 1528 203 1530 207
rect 1534 203 1537 207
rect 1542 203 1544 207
rect 1574 102 1577 1158
rect 1590 842 1593 928
rect 1598 912 1601 1198
rect 1598 862 1601 888
rect 1606 772 1609 1148
rect 1622 942 1625 968
rect 1582 742 1585 758
rect 1598 181 1601 748
rect 1614 662 1617 758
rect 1622 442 1625 848
rect 1630 822 1633 1218
rect 1646 1142 1649 1368
rect 1638 811 1641 1128
rect 1654 1072 1657 1328
rect 1662 1072 1665 1078
rect 1630 808 1641 811
rect 1646 1068 1654 1071
rect 1598 178 1606 181
rect 1630 142 1633 808
rect 1638 532 1641 728
rect 1646 662 1649 1068
rect 1646 562 1649 658
rect 1646 452 1649 558
rect 1646 372 1649 448
rect 1654 422 1657 938
rect 1662 852 1665 858
rect 1662 672 1665 678
rect 1638 112 1641 258
rect 1670 152 1673 1738
rect 1902 1672 1905 1718
rect 1694 1492 1697 1598
rect 1934 1562 1937 1758
rect 1966 1732 1969 1768
rect 1690 1268 1694 1271
rect 1710 1242 1713 1448
rect 1726 1408 1734 1411
rect 1726 1242 1729 1408
rect 1698 1078 1702 1081
rect 1718 1062 1721 1238
rect 1734 1212 1737 1398
rect 1742 1262 1745 1468
rect 1750 1132 1753 1528
rect 1826 1498 1833 1501
rect 1830 1452 1833 1498
rect 1794 1338 1798 1341
rect 1766 1291 1769 1298
rect 1762 1288 1769 1291
rect 1826 1288 1830 1291
rect 1838 1252 1841 1498
rect 1854 1442 1857 1458
rect 1902 1452 1905 1538
rect 1966 1512 1969 1728
rect 1890 1288 1894 1291
rect 1726 1082 1729 1088
rect 1802 1048 1809 1051
rect 1678 672 1681 678
rect 1686 662 1689 828
rect 1694 732 1697 988
rect 1762 868 1766 871
rect 1702 742 1705 868
rect 1806 722 1809 1048
rect 1886 552 1889 1218
rect 1902 422 1905 1448
rect 1958 1342 1961 1418
rect 1974 1342 1977 1638
rect 2014 1452 2017 1658
rect 1998 1412 2001 1428
rect 1910 1012 1913 1218
rect 1914 858 1918 861
rect 1926 502 1929 1058
rect 1934 732 1937 1098
rect 1942 752 1945 1118
rect 1950 662 1953 858
rect 1934 542 1937 658
rect 1958 462 1961 1338
rect 1862 418 1870 421
rect 1710 292 1713 418
rect 1718 262 1721 288
rect 1798 272 1801 298
rect 1862 252 1865 418
rect 1966 312 1969 1298
rect 1974 332 1977 1338
rect 1990 1301 1993 1358
rect 1986 1298 1993 1301
rect 1998 262 2001 1408
rect 2022 1282 2025 1378
rect 2022 1272 2025 1278
rect 2006 572 2009 1028
rect 2014 862 2017 868
rect 2014 682 2017 688
rect 2014 482 2017 658
rect 2022 472 2025 528
rect 1990 11 1993 198
rect 2030 12 2033 1368
rect 2046 1272 2049 1288
rect 2038 522 2041 1048
rect 2038 472 2041 488
rect 2046 62 2049 508
rect 1990 8 1998 11
rect 496 3 498 7
rect 502 3 505 7
rect 510 3 512 7
rect 1528 3 1530 7
rect 1534 3 1537 7
rect 1542 3 1544 7
<< m5contact >>
rect -18 1818 -14 1822
rect 498 1803 502 1807
rect 505 1803 506 1807
rect 506 1803 509 1807
rect 1530 1803 1534 1807
rect 1537 1803 1538 1807
rect 1538 1803 1541 1807
rect 22 1798 26 1802
rect 1018 1703 1022 1707
rect 1025 1703 1026 1707
rect 1026 1703 1029 1707
rect 182 668 186 672
rect 158 368 162 372
rect 318 1058 322 1062
rect 214 368 218 372
rect 174 258 178 262
rect 438 1288 442 1292
rect 430 1068 434 1072
rect 294 348 298 352
rect 498 1603 502 1607
rect 505 1603 506 1607
rect 506 1603 509 1607
rect 498 1403 502 1407
rect 505 1403 506 1407
rect 506 1403 509 1407
rect 494 1288 498 1292
rect 470 1258 474 1262
rect 498 1203 502 1207
rect 505 1203 506 1207
rect 506 1203 509 1207
rect 478 948 482 952
rect 498 1003 502 1007
rect 505 1003 506 1007
rect 506 1003 509 1007
rect 498 803 502 807
rect 505 803 506 807
rect 506 803 509 807
rect 590 1268 594 1272
rect 502 758 506 762
rect 498 603 502 607
rect 505 603 506 607
rect 506 603 509 607
rect 382 358 386 362
rect 406 348 410 352
rect 498 403 502 407
rect 505 403 506 407
rect 506 403 509 407
rect 486 338 490 342
rect 566 728 570 732
rect 590 938 594 942
rect 662 1288 666 1292
rect 638 928 642 932
rect 566 438 570 442
rect 630 668 634 672
rect 638 538 642 542
rect 614 358 618 362
rect 686 1008 690 1012
rect 550 258 554 262
rect 502 248 506 252
rect 606 248 610 252
rect 498 203 502 207
rect 505 203 506 207
rect 506 203 509 207
rect 718 758 722 762
rect 758 948 762 952
rect 718 748 722 752
rect 750 748 754 752
rect 742 738 746 742
rect 1018 1503 1022 1507
rect 1025 1503 1026 1507
rect 1026 1503 1029 1507
rect 814 1318 818 1322
rect 838 1278 842 1282
rect 862 1278 866 1282
rect 894 1278 898 1282
rect 782 848 786 852
rect 766 748 770 752
rect 782 738 786 742
rect 774 728 778 732
rect 774 718 778 722
rect 702 298 706 302
rect 726 268 730 272
rect 774 258 778 262
rect 822 738 826 742
rect 846 668 850 672
rect 878 748 882 752
rect 870 518 874 522
rect 814 368 818 372
rect 822 278 826 282
rect 886 458 890 462
rect 934 1068 938 1072
rect 990 1318 994 1322
rect 934 938 938 942
rect 910 728 914 732
rect 902 718 906 722
rect 926 658 930 662
rect 998 868 1002 872
rect 1018 1303 1022 1307
rect 1025 1303 1026 1307
rect 1026 1303 1029 1307
rect 1018 1103 1022 1107
rect 1025 1103 1026 1107
rect 1026 1103 1029 1107
rect 1018 903 1022 907
rect 1025 903 1026 907
rect 1026 903 1029 907
rect 910 488 914 492
rect 998 688 1002 692
rect 918 278 922 282
rect 942 278 946 282
rect 974 468 978 472
rect 958 338 962 342
rect 1018 703 1022 707
rect 1025 703 1026 707
rect 1026 703 1029 707
rect 1062 1258 1066 1262
rect 1046 1008 1050 1012
rect 1054 868 1058 872
rect 1018 503 1022 507
rect 1025 503 1026 507
rect 1026 503 1029 507
rect 1062 738 1066 742
rect 1046 468 1050 472
rect 1018 303 1022 307
rect 1025 303 1026 307
rect 1026 303 1029 307
rect 1006 298 1010 302
rect 926 258 930 262
rect 1046 458 1050 462
rect 1054 338 1058 342
rect 1046 288 1050 292
rect 1094 1278 1098 1282
rect 1530 1603 1534 1607
rect 1537 1603 1538 1607
rect 1538 1603 1541 1607
rect 1222 1348 1226 1352
rect 1182 1138 1186 1142
rect 1078 498 1082 502
rect 1094 498 1098 502
rect 1086 478 1090 482
rect 1094 368 1098 372
rect 1150 518 1154 522
rect 1134 488 1138 492
rect 1126 368 1130 372
rect 1166 338 1170 342
rect 1174 268 1178 272
rect 1206 538 1210 542
rect 1018 103 1022 107
rect 1025 103 1026 107
rect 1026 103 1029 107
rect 1366 1348 1370 1352
rect 1358 1298 1362 1302
rect 1302 1138 1306 1142
rect 1390 868 1394 872
rect 1286 678 1290 682
rect 1342 678 1346 682
rect 1358 658 1362 662
rect 1530 1403 1534 1407
rect 1537 1403 1538 1407
rect 1538 1403 1541 1407
rect 1518 1298 1522 1302
rect 1446 858 1450 862
rect 1422 738 1426 742
rect 1446 738 1450 742
rect 1438 728 1442 732
rect 1462 678 1466 682
rect 1550 1288 1554 1292
rect 1582 1268 1586 1272
rect 1530 1203 1534 1207
rect 1537 1203 1538 1207
rect 1538 1203 1541 1207
rect 1530 1003 1534 1007
rect 1537 1003 1538 1007
rect 1538 1003 1541 1007
rect 1534 928 1538 932
rect 1530 803 1534 807
rect 1537 803 1538 807
rect 1538 803 1541 807
rect 1550 738 1554 742
rect 1486 488 1490 492
rect 1530 603 1534 607
rect 1537 603 1538 607
rect 1538 603 1541 607
rect 1246 258 1250 262
rect 1566 438 1570 442
rect 1530 403 1534 407
rect 1537 403 1538 407
rect 1538 403 1541 407
rect 1530 203 1534 207
rect 1537 203 1538 207
rect 1538 203 1541 207
rect 1598 858 1602 862
rect 1582 738 1586 742
rect 1662 1068 1666 1072
rect 1662 858 1666 862
rect 1662 678 1666 682
rect 1694 1268 1698 1272
rect 1694 1078 1698 1082
rect 1798 1338 1802 1342
rect 1766 1298 1770 1302
rect 1830 1288 1834 1292
rect 1886 1288 1890 1292
rect 1726 1078 1730 1082
rect 1678 668 1682 672
rect 1758 868 1762 872
rect 1958 1338 1962 1342
rect 1918 858 1922 862
rect 1718 258 1722 262
rect 2022 1268 2026 1272
rect 2014 868 2018 872
rect 2014 688 2018 692
rect 498 3 502 7
rect 505 3 506 7
rect 506 3 509 7
rect 1530 3 1534 7
rect 1537 3 1538 7
rect 1538 3 1541 7
<< metal5 >>
rect -26 1818 -18 1821
rect -26 1801 -23 1818
rect 502 1803 505 1807
rect 501 1802 506 1803
rect 511 1802 512 1807
rect 1534 1803 1537 1807
rect 1533 1802 1538 1803
rect 1543 1802 1544 1807
rect -26 1798 22 1801
rect 1022 1703 1025 1707
rect 1021 1702 1026 1703
rect 1031 1702 1032 1707
rect 502 1603 505 1607
rect 501 1602 506 1603
rect 511 1602 512 1607
rect 1534 1603 1537 1607
rect 1533 1602 1538 1603
rect 1543 1602 1544 1607
rect 1022 1503 1025 1507
rect 1021 1502 1026 1503
rect 1031 1502 1032 1507
rect 502 1403 505 1407
rect 501 1402 506 1403
rect 511 1402 512 1407
rect 1534 1403 1537 1407
rect 1533 1402 1538 1403
rect 1543 1402 1544 1407
rect 1226 1348 1366 1351
rect 1802 1338 1958 1341
rect 818 1318 990 1321
rect 1022 1303 1025 1307
rect 1021 1302 1026 1303
rect 1031 1302 1032 1307
rect 1362 1298 1518 1301
rect 1522 1298 1766 1301
rect 442 1288 494 1291
rect 666 1288 1550 1291
rect 1834 1288 1886 1291
rect 842 1278 862 1281
rect 898 1278 1094 1281
rect 594 1268 1582 1271
rect 1698 1268 2022 1271
rect 474 1258 1062 1261
rect 502 1203 505 1207
rect 501 1202 506 1203
rect 511 1202 512 1207
rect 1534 1203 1537 1207
rect 1533 1202 1538 1203
rect 1543 1202 1544 1207
rect 1186 1138 1302 1141
rect 1022 1103 1025 1107
rect 1021 1102 1026 1103
rect 1031 1102 1032 1107
rect 1698 1078 1726 1081
rect 938 1068 1662 1071
rect 430 1061 433 1068
rect 322 1058 433 1061
rect 690 1008 1046 1011
rect 502 1003 505 1007
rect 501 1002 506 1003
rect 511 1002 512 1007
rect 1534 1003 1537 1007
rect 1533 1002 1538 1003
rect 1543 1002 1544 1007
rect 482 948 758 951
rect 594 938 934 941
rect 642 928 1534 931
rect 1022 903 1025 907
rect 1021 902 1026 903
rect 1031 902 1032 907
rect 1002 868 1054 871
rect 1394 868 1758 871
rect 1450 858 1598 861
rect 2014 861 2017 868
rect 1922 858 2017 861
rect 1662 851 1665 858
rect 786 848 1665 851
rect 502 803 505 807
rect 501 802 506 803
rect 511 802 512 807
rect 1534 803 1537 807
rect 1533 802 1538 803
rect 1543 802 1544 807
rect 506 758 718 761
rect 722 748 750 751
rect 770 748 878 751
rect 746 738 782 741
rect 826 738 1062 741
rect 1426 738 1446 741
rect 1554 738 1582 741
rect 570 728 774 731
rect 914 728 1438 731
rect 778 718 902 721
rect 1022 703 1025 707
rect 1021 702 1026 703
rect 1031 702 1032 707
rect 1002 688 2014 691
rect 1290 678 1342 681
rect 1466 678 1662 681
rect 186 668 630 671
rect 850 668 1678 671
rect 930 658 1358 661
rect 502 603 505 607
rect 501 602 506 603
rect 511 602 512 607
rect 1534 603 1537 607
rect 1533 602 1538 603
rect 1543 602 1544 607
rect 642 538 1206 541
rect 874 518 1150 521
rect 1022 503 1025 507
rect 1021 502 1026 503
rect 1031 502 1032 507
rect 1082 498 1094 501
rect 914 488 1134 491
rect 1486 481 1489 488
rect 1090 478 1489 481
rect 978 468 1046 471
rect 890 458 1046 461
rect 570 438 1566 441
rect 502 403 505 407
rect 501 402 506 403
rect 511 402 512 407
rect 1534 403 1537 407
rect 1533 402 1538 403
rect 1543 402 1544 407
rect 162 368 214 371
rect 218 368 814 371
rect 1098 368 1126 371
rect 386 358 614 361
rect 298 348 406 351
rect 490 338 958 341
rect 1058 338 1166 341
rect 1022 303 1025 307
rect 1021 302 1026 303
rect 1031 302 1032 307
rect 706 298 1006 301
rect 826 278 918 281
rect 1046 281 1049 288
rect 946 278 1049 281
rect 730 268 1174 271
rect 178 258 550 261
rect 778 258 926 261
rect 1250 258 1718 261
rect 506 248 606 251
rect 502 203 505 207
rect 501 202 506 203
rect 511 202 512 207
rect 1534 203 1537 207
rect 1533 202 1538 203
rect 1543 202 1544 207
rect 1022 103 1025 107
rect 1021 102 1026 103
rect 1031 102 1032 107
rect 502 3 505 7
rect 501 2 506 3
rect 511 2 512 7
rect 1534 3 1537 7
rect 1533 2 1538 3
rect 1543 2 1544 7
<< m6contact >>
rect 496 1803 498 1807
rect 498 1803 501 1807
rect 506 1803 509 1807
rect 509 1803 511 1807
rect 496 1802 501 1803
rect 506 1802 511 1803
rect 1528 1803 1530 1807
rect 1530 1803 1533 1807
rect 1538 1803 1541 1807
rect 1541 1803 1543 1807
rect 1528 1802 1533 1803
rect 1538 1802 1543 1803
rect 1016 1703 1018 1707
rect 1018 1703 1021 1707
rect 1026 1703 1029 1707
rect 1029 1703 1031 1707
rect 1016 1702 1021 1703
rect 1026 1702 1031 1703
rect 496 1603 498 1607
rect 498 1603 501 1607
rect 506 1603 509 1607
rect 509 1603 511 1607
rect 496 1602 501 1603
rect 506 1602 511 1603
rect 1528 1603 1530 1607
rect 1530 1603 1533 1607
rect 1538 1603 1541 1607
rect 1541 1603 1543 1607
rect 1528 1602 1533 1603
rect 1538 1602 1543 1603
rect 1016 1503 1018 1507
rect 1018 1503 1021 1507
rect 1026 1503 1029 1507
rect 1029 1503 1031 1507
rect 1016 1502 1021 1503
rect 1026 1502 1031 1503
rect 496 1403 498 1407
rect 498 1403 501 1407
rect 506 1403 509 1407
rect 509 1403 511 1407
rect 496 1402 501 1403
rect 506 1402 511 1403
rect 1528 1403 1530 1407
rect 1530 1403 1533 1407
rect 1538 1403 1541 1407
rect 1541 1403 1543 1407
rect 1528 1402 1533 1403
rect 1538 1402 1543 1403
rect 1016 1303 1018 1307
rect 1018 1303 1021 1307
rect 1026 1303 1029 1307
rect 1029 1303 1031 1307
rect 1016 1302 1021 1303
rect 1026 1302 1031 1303
rect 496 1203 498 1207
rect 498 1203 501 1207
rect 506 1203 509 1207
rect 509 1203 511 1207
rect 496 1202 501 1203
rect 506 1202 511 1203
rect 1528 1203 1530 1207
rect 1530 1203 1533 1207
rect 1538 1203 1541 1207
rect 1541 1203 1543 1207
rect 1528 1202 1533 1203
rect 1538 1202 1543 1203
rect 1016 1103 1018 1107
rect 1018 1103 1021 1107
rect 1026 1103 1029 1107
rect 1029 1103 1031 1107
rect 1016 1102 1021 1103
rect 1026 1102 1031 1103
rect 496 1003 498 1007
rect 498 1003 501 1007
rect 506 1003 509 1007
rect 509 1003 511 1007
rect 496 1002 501 1003
rect 506 1002 511 1003
rect 1528 1003 1530 1007
rect 1530 1003 1533 1007
rect 1538 1003 1541 1007
rect 1541 1003 1543 1007
rect 1528 1002 1533 1003
rect 1538 1002 1543 1003
rect 1016 903 1018 907
rect 1018 903 1021 907
rect 1026 903 1029 907
rect 1029 903 1031 907
rect 1016 902 1021 903
rect 1026 902 1031 903
rect 496 803 498 807
rect 498 803 501 807
rect 506 803 509 807
rect 509 803 511 807
rect 496 802 501 803
rect 506 802 511 803
rect 1528 803 1530 807
rect 1530 803 1533 807
rect 1538 803 1541 807
rect 1541 803 1543 807
rect 1528 802 1533 803
rect 1538 802 1543 803
rect 1016 703 1018 707
rect 1018 703 1021 707
rect 1026 703 1029 707
rect 1029 703 1031 707
rect 1016 702 1021 703
rect 1026 702 1031 703
rect 496 603 498 607
rect 498 603 501 607
rect 506 603 509 607
rect 509 603 511 607
rect 496 602 501 603
rect 506 602 511 603
rect 1528 603 1530 607
rect 1530 603 1533 607
rect 1538 603 1541 607
rect 1541 603 1543 607
rect 1528 602 1533 603
rect 1538 602 1543 603
rect 1016 503 1018 507
rect 1018 503 1021 507
rect 1026 503 1029 507
rect 1029 503 1031 507
rect 1016 502 1021 503
rect 1026 502 1031 503
rect 496 403 498 407
rect 498 403 501 407
rect 506 403 509 407
rect 509 403 511 407
rect 496 402 501 403
rect 506 402 511 403
rect 1528 403 1530 407
rect 1530 403 1533 407
rect 1538 403 1541 407
rect 1541 403 1543 407
rect 1528 402 1533 403
rect 1538 402 1543 403
rect 1016 303 1018 307
rect 1018 303 1021 307
rect 1026 303 1029 307
rect 1029 303 1031 307
rect 1016 302 1021 303
rect 1026 302 1031 303
rect 496 203 498 207
rect 498 203 501 207
rect 506 203 509 207
rect 509 203 511 207
rect 496 202 501 203
rect 506 202 511 203
rect 1528 203 1530 207
rect 1530 203 1533 207
rect 1538 203 1541 207
rect 1541 203 1543 207
rect 1528 202 1533 203
rect 1538 202 1543 203
rect 1016 103 1018 107
rect 1018 103 1021 107
rect 1026 103 1029 107
rect 1029 103 1031 107
rect 1016 102 1021 103
rect 1026 102 1031 103
rect 496 3 498 7
rect 498 3 501 7
rect 506 3 509 7
rect 509 3 511 7
rect 496 2 501 3
rect 506 2 511 3
rect 1528 3 1530 7
rect 1530 3 1533 7
rect 1538 3 1541 7
rect 1541 3 1543 7
rect 1528 2 1533 3
rect 1538 2 1543 3
<< metal6 >>
rect 496 1807 512 1830
rect 501 1802 506 1807
rect 511 1802 512 1807
rect 496 1607 512 1802
rect 501 1602 506 1607
rect 511 1602 512 1607
rect 496 1407 512 1602
rect 501 1402 506 1407
rect 511 1402 512 1407
rect 496 1207 512 1402
rect 501 1202 506 1207
rect 511 1202 512 1207
rect 496 1007 512 1202
rect 501 1002 506 1007
rect 511 1002 512 1007
rect 496 807 512 1002
rect 501 802 506 807
rect 511 802 512 807
rect 496 607 512 802
rect 501 602 506 607
rect 511 602 512 607
rect 496 407 512 602
rect 501 402 506 407
rect 511 402 512 407
rect 496 207 512 402
rect 501 202 506 207
rect 511 202 512 207
rect 496 7 512 202
rect 501 2 506 7
rect 511 2 512 7
rect 496 -30 512 2
rect 1016 1707 1032 1830
rect 1021 1702 1026 1707
rect 1031 1702 1032 1707
rect 1016 1507 1032 1702
rect 1021 1502 1026 1507
rect 1031 1502 1032 1507
rect 1016 1307 1032 1502
rect 1021 1302 1026 1307
rect 1031 1302 1032 1307
rect 1016 1107 1032 1302
rect 1021 1102 1026 1107
rect 1031 1102 1032 1107
rect 1016 907 1032 1102
rect 1021 902 1026 907
rect 1031 902 1032 907
rect 1016 707 1032 902
rect 1021 702 1026 707
rect 1031 702 1032 707
rect 1016 507 1032 702
rect 1021 502 1026 507
rect 1031 502 1032 507
rect 1016 307 1032 502
rect 1021 302 1026 307
rect 1031 302 1032 307
rect 1016 107 1032 302
rect 1021 102 1026 107
rect 1031 102 1032 107
rect 1016 -30 1032 102
rect 1528 1807 1544 1830
rect 1533 1802 1538 1807
rect 1543 1802 1544 1807
rect 1528 1607 1544 1802
rect 1533 1602 1538 1607
rect 1543 1602 1544 1607
rect 1528 1407 1544 1602
rect 1533 1402 1538 1407
rect 1543 1402 1544 1407
rect 1528 1207 1544 1402
rect 1533 1202 1538 1207
rect 1543 1202 1544 1207
rect 1528 1007 1544 1202
rect 1533 1002 1538 1007
rect 1543 1002 1544 1007
rect 1528 807 1544 1002
rect 1533 802 1538 807
rect 1543 802 1544 807
rect 1528 607 1544 802
rect 1533 602 1538 607
rect 1543 602 1544 607
rect 1528 407 1544 602
rect 1533 402 1538 407
rect 1543 402 1544 407
rect 1528 207 1544 402
rect 1533 202 1538 207
rect 1543 202 1544 207
rect 1528 7 1544 202
rect 1533 2 1538 7
rect 1543 2 1544 7
rect 1528 -30 1544 2
use CLKBUF1  CLKBUF1_9
timestamp 1713260442
transform 1 0 4 0 -1 105
box -2 -3 74 103
use CLKBUF1  CLKBUF1_5
timestamp 1713260442
transform 1 0 76 0 -1 105
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_42
timestamp 1713260442
transform 1 0 148 0 -1 105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_24
timestamp 1713260442
transform 1 0 4 0 1 105
box -2 -3 98 103
use AOI21X1  AOI21X1_91
timestamp 1713260442
transform 1 0 100 0 1 105
box -2 -3 34 103
use NOR2X1  NOR2X1_65
timestamp 1713260442
transform -1 0 156 0 1 105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_115
timestamp 1713260442
transform 1 0 156 0 1 105
box -2 -3 98 103
use NOR2X1  NOR2X1_14
timestamp 1713260442
transform 1 0 244 0 -1 105
box -2 -3 26 103
use AOI21X1  AOI21X1_11
timestamp 1713260442
transform -1 0 300 0 -1 105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_3
timestamp 1713260442
transform 1 0 300 0 -1 105
box -2 -3 98 103
use OAI21X1  OAI21X1_19
timestamp 1713260442
transform 1 0 252 0 1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_22
timestamp 1713260442
transform -1 0 308 0 1 105
box -2 -3 26 103
use OAI21X1  OAI21X1_160
timestamp 1713260442
transform 1 0 308 0 1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_92
timestamp 1713260442
transform -1 0 364 0 1 105
box -2 -3 26 103
use INVX1  INVX1_34
timestamp 1713260442
transform 1 0 364 0 1 105
box -2 -3 18 103
use NAND2X1  NAND2X1_5
timestamp 1713260442
transform 1 0 380 0 1 105
box -2 -3 26 103
use OAI21X1  OAI21X1_5
timestamp 1713260442
transform -1 0 428 0 -1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_47
timestamp 1713260442
transform 1 0 516 0 1 105
box -2 -3 34 103
use FILL  FILL_1_0_1
timestamp 1713260442
transform 1 0 508 0 1 105
box -2 -3 10 103
use FILL  FILL_1_0_0
timestamp 1713260442
transform 1 0 500 0 1 105
box -2 -3 10 103
use FILL  FILL_0_0_1
timestamp 1713260442
transform 1 0 532 0 -1 105
box -2 -3 10 103
use FILL  FILL_0_0_0
timestamp 1713260442
transform 1 0 524 0 -1 105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_87
timestamp 1713260442
transform 1 0 404 0 1 105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_122
timestamp 1713260442
transform 1 0 540 0 -1 105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_37
timestamp 1713260442
transform -1 0 524 0 -1 105
box -2 -3 98 103
use NAND2X1  NAND2X1_13
timestamp 1713260442
transform 1 0 636 0 -1 105
box -2 -3 26 103
use OAI21X1  OAI21X1_10
timestamp 1713260442
transform -1 0 692 0 -1 105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_128
timestamp 1713260442
transform 1 0 692 0 -1 105
box -2 -3 98 103
use NAND2X1  NAND2X1_50
timestamp 1713260442
transform -1 0 572 0 1 105
box -2 -3 26 103
use NOR2X1  NOR2X1_41
timestamp 1713260442
transform 1 0 572 0 1 105
box -2 -3 26 103
use NOR2X1  NOR2X1_39
timestamp 1713260442
transform -1 0 620 0 1 105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_59
timestamp 1713260442
transform -1 0 716 0 1 105
box -2 -3 98 103
use OAI21X1  OAI21X1_16
timestamp 1713260442
transform 1 0 716 0 1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_19
timestamp 1713260442
transform -1 0 812 0 -1 105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_101
timestamp 1713260442
transform -1 0 908 0 -1 105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_117
timestamp 1713260442
transform -1 0 1004 0 -1 105
box -2 -3 98 103
use OAI21X1  OAI21X1_80
timestamp 1713260442
transform 1 0 748 0 1 105
box -2 -3 34 103
use OAI22X1  OAI22X1_1
timestamp 1713260442
transform -1 0 820 0 1 105
box -2 -3 42 103
use INVX1  INVX1_36
timestamp 1713260442
transform 1 0 820 0 1 105
box -2 -3 18 103
use NAND2X1  NAND2X1_24
timestamp 1713260442
transform 1 0 836 0 1 105
box -2 -3 26 103
use OAI21X1  OAI21X1_21
timestamp 1713260442
transform -1 0 892 0 1 105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_100
timestamp 1713260442
transform 1 0 892 0 1 105
box -2 -3 98 103
use FILL  FILL_0_1_0
timestamp 1713260442
transform -1 0 1012 0 -1 105
box -2 -3 10 103
use FILL  FILL_0_1_1
timestamp 1713260442
transform -1 0 1020 0 -1 105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_123
timestamp 1713260442
transform -1 0 1116 0 -1 105
box -2 -3 98 103
use INVX1  INVX1_30
timestamp 1713260442
transform -1 0 1004 0 1 105
box -2 -3 18 103
use NOR2X1  NOR2X1_38
timestamp 1713260442
transform 1 0 1004 0 1 105
box -2 -3 26 103
use FILL  FILL_1_1_0
timestamp 1713260442
transform -1 0 1036 0 1 105
box -2 -3 10 103
use FILL  FILL_1_1_1
timestamp 1713260442
transform -1 0 1044 0 1 105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_21
timestamp 1713260442
transform -1 0 1140 0 1 105
box -2 -3 98 103
use NAND2X1  NAND2X1_14
timestamp 1713260442
transform 1 0 1116 0 -1 105
box -2 -3 26 103
use OAI21X1  OAI21X1_11
timestamp 1713260442
transform -1 0 1172 0 -1 105
box -2 -3 34 103
use NOR2X1  NOR2X1_15
timestamp 1713260442
transform -1 0 1196 0 -1 105
box -2 -3 26 103
use AOI21X1  AOI21X1_12
timestamp 1713260442
transform -1 0 1228 0 -1 105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_43
timestamp 1713260442
transform -1 0 1324 0 -1 105
box -2 -3 98 103
use NAND2X1  NAND2X1_96
timestamp 1713260442
transform 1 0 1140 0 1 105
box -2 -3 26 103
use OAI21X1  OAI21X1_164
timestamp 1713260442
transform -1 0 1196 0 1 105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_7
timestamp 1713260442
transform 1 0 1196 0 1 105
box -2 -3 98 103
use INVX1  INVX1_18
timestamp 1713260442
transform -1 0 1340 0 -1 105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_50
timestamp 1713260442
transform -1 0 1436 0 -1 105
box -2 -3 98 103
use CLKBUF1  CLKBUF1_12
timestamp 1713260442
transform 1 0 1436 0 -1 105
box -2 -3 74 103
use CLKBUF1  CLKBUF1_11
timestamp 1713260442
transform -1 0 1364 0 1 105
box -2 -3 74 103
use MUX2X1  MUX2X1_2
timestamp 1713260442
transform 1 0 1364 0 1 105
box -2 -3 50 103
use NOR2X1  NOR2X1_5
timestamp 1713260442
transform 1 0 1412 0 1 105
box -2 -3 26 103
use AOI21X1  AOI21X1_3
timestamp 1713260442
transform -1 0 1468 0 1 105
box -2 -3 34 103
use FILL  FILL_0_2_0
timestamp 1713260442
transform -1 0 1516 0 -1 105
box -2 -3 10 103
use FILL  FILL_0_2_1
timestamp 1713260442
transform -1 0 1524 0 -1 105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_75
timestamp 1713260442
transform -1 0 1620 0 -1 105
box -2 -3 98 103
use INVX1  INVX1_5
timestamp 1713260442
transform 1 0 1620 0 -1 105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_74
timestamp 1713260442
transform -1 0 1564 0 1 105
box -2 -3 98 103
use FILL  FILL_1_2_0
timestamp 1713260442
transform 1 0 1564 0 1 105
box -2 -3 10 103
use FILL  FILL_1_2_1
timestamp 1713260442
transform 1 0 1572 0 1 105
box -2 -3 10 103
use NOR2X1  NOR2X1_6
timestamp 1713260442
transform 1 0 1580 0 1 105
box -2 -3 26 103
use AOI21X1  AOI21X1_4
timestamp 1713260442
transform -1 0 1636 0 1 105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_51
timestamp 1713260442
transform -1 0 1732 0 -1 105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_73
timestamp 1713260442
transform -1 0 1828 0 -1 105
box -2 -3 98 103
use NOR2X1  NOR2X1_1
timestamp 1713260442
transform 1 0 1636 0 1 105
box -2 -3 26 103
use AOI21X1  AOI21X1_1
timestamp 1713260442
transform -1 0 1692 0 1 105
box -2 -3 34 103
use CLKBUF1  CLKBUF1_10
timestamp 1713260442
transform 1 0 1692 0 1 105
box -2 -3 74 103
use NOR2X1  NOR2X1_4
timestamp 1713260442
transform 1 0 1764 0 1 105
box -2 -3 26 103
use AOI21X1  AOI21X1_2
timestamp 1713260442
transform -1 0 1820 0 1 105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_11
timestamp 1713260442
transform -1 0 1924 0 -1 105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_49
timestamp 1713260442
transform 1 0 1924 0 -1 105
box -2 -3 98 103
use NOR2X1  NOR2X1_76
timestamp 1713260442
transform 1 0 1820 0 1 105
box -2 -3 26 103
use AOI21X1  AOI21X1_100
timestamp 1713260442
transform -1 0 1876 0 1 105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_25
timestamp 1713260442
transform 1 0 1876 0 1 105
box -2 -3 98 103
use BUFX2  BUFX2_13
timestamp 1713260442
transform 1 0 1972 0 1 105
box -2 -3 26 103
use INVX4  INVX4_1
timestamp 1713260442
transform 1 0 2020 0 -1 105
box -2 -3 26 103
use FILL  FILL_1_1
timestamp 1713260442
transform -1 0 2052 0 -1 105
box -2 -3 10 103
use INVX1  INVX1_10
timestamp 1713260442
transform -1 0 2012 0 1 105
box -2 -3 18 103
use BUFX2  BUFX2_12
timestamp 1713260442
transform 1 0 2012 0 1 105
box -2 -3 26 103
use FILL  FILL_2_1
timestamp 1713260442
transform 1 0 2036 0 1 105
box -2 -3 10 103
use FILL  FILL_2_2
timestamp 1713260442
transform 1 0 2044 0 1 105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_104
timestamp 1713260442
transform -1 0 100 0 -1 305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_19
timestamp 1713260442
transform -1 0 196 0 -1 305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_83
timestamp 1713260442
transform 1 0 196 0 -1 305
box -2 -3 98 103
use NAND2X1  NAND2X1_46
timestamp 1713260442
transform 1 0 292 0 -1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_43
timestamp 1713260442
transform -1 0 348 0 -1 305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_35
timestamp 1713260442
transform 1 0 348 0 -1 305
box -2 -3 98 103
use OAI21X1  OAI21X1_3
timestamp 1713260442
transform 1 0 444 0 -1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_3
timestamp 1713260442
transform -1 0 500 0 -1 305
box -2 -3 26 103
use FILL  FILL_2_0_0
timestamp 1713260442
transform -1 0 508 0 -1 305
box -2 -3 10 103
use FILL  FILL_2_0_1
timestamp 1713260442
transform -1 0 516 0 -1 305
box -2 -3 10 103
use BUFX4  BUFX4_46
timestamp 1713260442
transform -1 0 548 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_143
timestamp 1713260442
transform 1 0 548 0 -1 305
box -2 -3 34 103
use AOI21X1  AOI21X1_81
timestamp 1713260442
transform -1 0 612 0 -1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_40
timestamp 1713260442
transform 1 0 612 0 -1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_86
timestamp 1713260442
transform -1 0 668 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_107
timestamp 1713260442
transform 1 0 668 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_88
timestamp 1713260442
transform -1 0 732 0 -1 305
box -2 -3 34 103
use MUX2X1  MUX2X1_13
timestamp 1713260442
transform -1 0 780 0 -1 305
box -2 -3 50 103
use NAND2X1  NAND2X1_78
timestamp 1713260442
transform 1 0 780 0 -1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_152
timestamp 1713260442
transform -1 0 836 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_110
timestamp 1713260442
transform 1 0 836 0 -1 305
box -2 -3 34 103
use MUX2X1  MUX2X1_26
timestamp 1713260442
transform 1 0 868 0 -1 305
box -2 -3 50 103
use OAI21X1  OAI21X1_85
timestamp 1713260442
transform 1 0 916 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_84
timestamp 1713260442
transform 1 0 948 0 -1 305
box -2 -3 34 103
use MUX2X1  MUX2X1_25
timestamp 1713260442
transform 1 0 980 0 -1 305
box -2 -3 50 103
use FILL  FILL_2_1_0
timestamp 1713260442
transform -1 0 1036 0 -1 305
box -2 -3 10 103
use FILL  FILL_2_1_1
timestamp 1713260442
transform -1 0 1044 0 -1 305
box -2 -3 10 103
use AOI21X1  AOI21X1_60
timestamp 1713260442
transform -1 0 1076 0 -1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_62
timestamp 1713260442
transform 1 0 1076 0 -1 305
box -2 -3 26 103
use AOI21X1  AOI21X1_88
timestamp 1713260442
transform -1 0 1132 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_89
timestamp 1713260442
transform -1 0 1164 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_83
timestamp 1713260442
transform -1 0 1196 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_81
timestamp 1713260442
transform -1 0 1228 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_87
timestamp 1713260442
transform 1 0 1228 0 -1 305
box -2 -3 34 103
use AOI21X1  AOI21X1_40
timestamp 1713260442
transform 1 0 1260 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_72
timestamp 1713260442
transform -1 0 1324 0 -1 305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_66
timestamp 1713260442
transform -1 0 1420 0 -1 305
box -2 -3 98 103
use NOR2X1  NOR2X1_42
timestamp 1713260442
transform 1 0 1420 0 -1 305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_26
timestamp 1713260442
transform -1 0 1540 0 -1 305
box -2 -3 98 103
use FILL  FILL_2_2_0
timestamp 1713260442
transform 1 0 1540 0 -1 305
box -2 -3 10 103
use FILL  FILL_2_2_1
timestamp 1713260442
transform 1 0 1548 0 -1 305
box -2 -3 10 103
use AOI21X1  AOI21X1_18
timestamp 1713260442
transform 1 0 1556 0 -1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_22
timestamp 1713260442
transform 1 0 1588 0 -1 305
box -2 -3 26 103
use AOI21X1  AOI21X1_36
timestamp 1713260442
transform -1 0 1644 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_70
timestamp 1713260442
transform -1 0 1676 0 -1 305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_65
timestamp 1713260442
transform -1 0 1772 0 -1 305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_67
timestamp 1713260442
transform -1 0 1868 0 -1 305
box -2 -3 98 103
use MUX2X1  MUX2X1_8
timestamp 1713260442
transform 1 0 1868 0 -1 305
box -2 -3 50 103
use INVX2  INVX2_1
timestamp 1713260442
transform -1 0 1932 0 -1 305
box -2 -3 18 103
use INVX1  INVX1_16
timestamp 1713260442
transform -1 0 1948 0 -1 305
box -2 -3 18 103
use MUX2X1  MUX2X1_1
timestamp 1713260442
transform 1 0 1948 0 -1 305
box -2 -3 50 103
use BUFX2  BUFX2_10
timestamp 1713260442
transform -1 0 2020 0 -1 305
box -2 -3 26 103
use BUFX2  BUFX2_14
timestamp 1713260442
transform 1 0 2020 0 -1 305
box -2 -3 26 103
use FILL  FILL_3_1
timestamp 1713260442
transform -1 0 2052 0 -1 305
box -2 -3 10 103
use INVX1  INVX1_54
timestamp 1713260442
transform 1 0 4 0 1 305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_107
timestamp 1713260442
transform 1 0 20 0 1 305
box -2 -3 98 103
use MUX2X1  MUX2X1_29
timestamp 1713260442
transform -1 0 164 0 1 305
box -2 -3 50 103
use INVX1  INVX1_25
timestamp 1713260442
transform 1 0 164 0 1 305
box -2 -3 18 103
use MUX2X1  MUX2X1_14
timestamp 1713260442
transform 1 0 180 0 1 305
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_58
timestamp 1713260442
transform 1 0 228 0 1 305
box -2 -3 98 103
use OAI21X1  OAI21X1_151
timestamp 1713260442
transform 1 0 324 0 1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_76
timestamp 1713260442
transform 1 0 356 0 1 305
box -2 -3 26 103
use INVX1  INVX1_26
timestamp 1713260442
transform 1 0 380 0 1 305
box -2 -3 18 103
use AOI21X1  AOI21X1_48
timestamp 1713260442
transform 1 0 396 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_91
timestamp 1713260442
transform 1 0 428 0 1 305
box -2 -3 34 103
use AOI21X1  AOI21X1_49
timestamp 1713260442
transform 1 0 460 0 1 305
box -2 -3 34 103
use FILL  FILL_3_0_0
timestamp 1713260442
transform 1 0 492 0 1 305
box -2 -3 10 103
use FILL  FILL_3_0_1
timestamp 1713260442
transform 1 0 500 0 1 305
box -2 -3 10 103
use AOI21X1  AOI21X1_42
timestamp 1713260442
transform 1 0 508 0 1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_45
timestamp 1713260442
transform 1 0 540 0 1 305
box -2 -3 26 103
use NOR2X1  NOR2X1_53
timestamp 1713260442
transform 1 0 564 0 1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_75
timestamp 1713260442
transform -1 0 620 0 1 305
box -2 -3 34 103
use BUFX4  BUFX4_25
timestamp 1713260442
transform -1 0 652 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_153
timestamp 1713260442
transform 1 0 652 0 1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_80
timestamp 1713260442
transform -1 0 708 0 1 305
box -2 -3 26 103
use BUFX4  BUFX4_33
timestamp 1713260442
transform -1 0 740 0 1 305
box -2 -3 34 103
use INVX8  INVX8_2
timestamp 1713260442
transform -1 0 780 0 1 305
box -2 -3 42 103
use NOR2X1  NOR2X1_55
timestamp 1713260442
transform 1 0 780 0 1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_99
timestamp 1713260442
transform -1 0 836 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_157
timestamp 1713260442
transform 1 0 836 0 1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_87
timestamp 1713260442
transform -1 0 892 0 1 305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_64
timestamp 1713260442
transform -1 0 988 0 1 305
box -2 -3 98 103
use NOR2X1  NOR2X1_43
timestamp 1713260442
transform -1 0 1012 0 1 305
box -2 -3 26 103
use FILL  FILL_3_1_0
timestamp 1713260442
transform 1 0 1012 0 1 305
box -2 -3 10 103
use FILL  FILL_3_1_1
timestamp 1713260442
transform 1 0 1020 0 1 305
box -2 -3 10 103
use OAI22X1  OAI22X1_3
timestamp 1713260442
transform 1 0 1028 0 1 305
box -2 -3 42 103
use MUX2X1  MUX2X1_24
timestamp 1713260442
transform -1 0 1116 0 1 305
box -2 -3 50 103
use AOI21X1  AOI21X1_47
timestamp 1713260442
transform 1 0 1116 0 1 305
box -2 -3 34 103
use INVX1  INVX1_24
timestamp 1713260442
transform -1 0 1164 0 1 305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_99
timestamp 1713260442
transform -1 0 1260 0 1 305
box -2 -3 98 103
use NOR2X1  NOR2X1_68
timestamp 1713260442
transform 1 0 1260 0 1 305
box -2 -3 26 103
use AOI21X1  AOI21X1_93
timestamp 1713260442
transform -1 0 1316 0 1 305
box -2 -3 34 103
use MUX2X1  MUX2X1_16
timestamp 1713260442
transform -1 0 1364 0 1 305
box -2 -3 50 103
use INVX1  INVX1_20
timestamp 1713260442
transform -1 0 1380 0 1 305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_10
timestamp 1713260442
transform -1 0 1476 0 1 305
box -2 -3 98 103
use CLKBUF1  CLKBUF1_1
timestamp 1713260442
transform -1 0 1548 0 1 305
box -2 -3 74 103
use FILL  FILL_3_2_0
timestamp 1713260442
transform -1 0 1556 0 1 305
box -2 -3 10 103
use FILL  FILL_3_2_1
timestamp 1713260442
transform -1 0 1564 0 1 305
box -2 -3 10 103
use INVX1  INVX1_53
timestamp 1713260442
transform -1 0 1580 0 1 305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_16
timestamp 1713260442
transform -1 0 1676 0 1 305
box -2 -3 98 103
use NOR2X1  NOR2X1_67
timestamp 1713260442
transform 1 0 1676 0 1 305
box -2 -3 26 103
use AOI21X1  AOI21X1_92
timestamp 1713260442
transform -1 0 1732 0 1 305
box -2 -3 34 103
use MUX2X1  MUX2X1_15
timestamp 1713260442
transform 1 0 1732 0 1 305
box -2 -3 50 103
use INVX1  INVX1_12
timestamp 1713260442
transform -1 0 1796 0 1 305
box -2 -3 18 103
use NOR2X1  NOR2X1_69
timestamp 1713260442
transform 1 0 1796 0 1 305
box -2 -3 26 103
use AOI21X1  AOI21X1_94
timestamp 1713260442
transform -1 0 1852 0 1 305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_9
timestamp 1713260442
transform -1 0 1948 0 1 305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_71
timestamp 1713260442
transform -1 0 2044 0 1 305
box -2 -3 98 103
use FILL  FILL_4_1
timestamp 1713260442
transform 1 0 2044 0 1 305
box -2 -3 10 103
use CLKBUF1  CLKBUF1_7
timestamp 1713260442
transform 1 0 4 0 -1 505
box -2 -3 74 103
use NOR2X1  NOR2X1_20
timestamp 1713260442
transform 1 0 76 0 -1 505
box -2 -3 26 103
use AOI21X1  AOI21X1_17
timestamp 1713260442
transform -1 0 132 0 -1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_30
timestamp 1713260442
transform 1 0 132 0 -1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_27
timestamp 1713260442
transform -1 0 188 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_35
timestamp 1713260442
transform 1 0 188 0 -1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_38
timestamp 1713260442
transform -1 0 244 0 -1 505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_91
timestamp 1713260442
transform 1 0 244 0 -1 505
box -2 -3 98 103
use OAI21X1  OAI21X1_159
timestamp 1713260442
transform 1 0 340 0 -1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_91
timestamp 1713260442
transform -1 0 396 0 -1 505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_2
timestamp 1713260442
transform 1 0 396 0 -1 505
box -2 -3 98 103
use FILL  FILL_4_0_0
timestamp 1713260442
transform 1 0 492 0 -1 505
box -2 -3 10 103
use FILL  FILL_4_0_1
timestamp 1713260442
transform 1 0 500 0 -1 505
box -2 -3 10 103
use OAI21X1  OAI21X1_92
timestamp 1713260442
transform 1 0 508 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_93
timestamp 1713260442
transform 1 0 540 0 -1 505
box -2 -3 34 103
use BUFX4  BUFX4_29
timestamp 1713260442
transform 1 0 572 0 -1 505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_60
timestamp 1713260442
transform 1 0 604 0 -1 505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_103
timestamp 1713260442
transform 1 0 700 0 -1 505
box -2 -3 98 103
use INVX1  INVX1_48
timestamp 1713260442
transform 1 0 796 0 -1 505
box -2 -3 18 103
use MUX2X1  MUX2X1_28
timestamp 1713260442
transform -1 0 860 0 -1 505
box -2 -3 50 103
use NOR2X1  NOR2X1_48
timestamp 1713260442
transform -1 0 884 0 -1 505
box -2 -3 26 103
use AOI21X1  AOI21X1_52
timestamp 1713260442
transform 1 0 884 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_132
timestamp 1713260442
transform 1 0 916 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_144
timestamp 1713260442
transform -1 0 980 0 -1 505
box -2 -3 34 103
use BUFX4  BUFX4_24
timestamp 1713260442
transform 1 0 980 0 -1 505
box -2 -3 34 103
use FILL  FILL_4_1_0
timestamp 1713260442
transform 1 0 1012 0 -1 505
box -2 -3 10 103
use FILL  FILL_4_1_1
timestamp 1713260442
transform 1 0 1020 0 -1 505
box -2 -3 10 103
use AOI21X1  AOI21X1_33
timestamp 1713260442
transform 1 0 1028 0 -1 505
box -2 -3 34 103
use AOI21X1  AOI21X1_80
timestamp 1713260442
transform 1 0 1060 0 -1 505
box -2 -3 34 103
use AOI21X1  AOI21X1_74
timestamp 1713260442
transform -1 0 1124 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_90
timestamp 1713260442
transform -1 0 1156 0 -1 505
box -2 -3 34 103
use NOR2X1  NOR2X1_64
timestamp 1713260442
transform -1 0 1180 0 -1 505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_23
timestamp 1713260442
transform -1 0 1276 0 -1 505
box -2 -3 98 103
use OAI21X1  OAI21X1_98
timestamp 1713260442
transform -1 0 1308 0 -1 505
box -2 -3 34 103
use BUFX4  BUFX4_26
timestamp 1713260442
transform -1 0 1340 0 -1 505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_27
timestamp 1713260442
transform -1 0 1436 0 -1 505
box -2 -3 98 103
use NOR2X1  NOR2X1_23
timestamp 1713260442
transform 1 0 1436 0 -1 505
box -2 -3 26 103
use AOI21X1  AOI21X1_19
timestamp 1713260442
transform -1 0 1492 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_142
timestamp 1713260442
transform -1 0 1524 0 -1 505
box -2 -3 34 103
use FILL  FILL_4_2_0
timestamp 1713260442
transform -1 0 1532 0 -1 505
box -2 -3 10 103
use FILL  FILL_4_2_1
timestamp 1713260442
transform -1 0 1540 0 -1 505
box -2 -3 10 103
use INVX4  INVX4_2
timestamp 1713260442
transform -1 0 1564 0 -1 505
box -2 -3 26 103
use MUX2X1  MUX2X1_21
timestamp 1713260442
transform 1 0 1564 0 -1 505
box -2 -3 50 103
use AOI21X1  AOI21X1_28
timestamp 1713260442
transform 1 0 1612 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_62
timestamp 1713260442
transform -1 0 1676 0 -1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_75
timestamp 1713260442
transform 1 0 1676 0 -1 505
box -2 -3 26 103
use NAND2X1  NAND2X1_77
timestamp 1713260442
transform -1 0 1724 0 -1 505
box -2 -3 26 103
use INVX4  INVX4_3
timestamp 1713260442
transform 1 0 1724 0 -1 505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_56
timestamp 1713260442
transform 1 0 1748 0 -1 505
box -2 -3 98 103
use INVX1  INVX1_51
timestamp 1713260442
transform 1 0 1844 0 -1 505
box -2 -3 18 103
use MUX2X1  MUX2X1_7
timestamp 1713260442
transform 1 0 1860 0 -1 505
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_72
timestamp 1713260442
transform 1 0 1908 0 -1 505
box -2 -3 98 103
use INVX4  INVX4_5
timestamp 1713260442
transform 1 0 2004 0 -1 505
box -2 -3 26 103
use NOR2X1  NOR2X1_73
timestamp 1713260442
transform 1 0 2028 0 -1 505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_48
timestamp 1713260442
transform 1 0 4 0 1 505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_93
timestamp 1713260442
transform 1 0 100 0 1 505
box -2 -3 98 103
use OAI21X1  OAI21X1_37
timestamp 1713260442
transform 1 0 196 0 1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_40
timestamp 1713260442
transform -1 0 252 0 1 505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_88
timestamp 1713260442
transform 1 0 252 0 1 505
box -2 -3 98 103
use NAND2X1  NAND2X1_52
timestamp 1713260442
transform 1 0 348 0 1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_48
timestamp 1713260442
transform -1 0 404 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_115
timestamp 1713260442
transform 1 0 404 0 1 505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_119
timestamp 1713260442
transform 1 0 436 0 1 505
box -2 -3 98 103
use FILL  FILL_5_0_0
timestamp 1713260442
transform 1 0 532 0 1 505
box -2 -3 10 103
use FILL  FILL_5_0_1
timestamp 1713260442
transform 1 0 540 0 1 505
box -2 -3 10 103
use OAI21X1  OAI21X1_23
timestamp 1713260442
transform 1 0 548 0 1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_26
timestamp 1713260442
transform -1 0 604 0 1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_74
timestamp 1713260442
transform -1 0 636 0 1 505
box -2 -3 34 103
use AOI21X1  AOI21X1_41
timestamp 1713260442
transform 1 0 636 0 1 505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_92
timestamp 1713260442
transform 1 0 668 0 1 505
box -2 -3 98 103
use OAI21X1  OAI21X1_36
timestamp 1713260442
transform 1 0 764 0 1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_39
timestamp 1713260442
transform -1 0 820 0 1 505
box -2 -3 26 103
use AOI21X1  AOI21X1_53
timestamp 1713260442
transform -1 0 852 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_100
timestamp 1713260442
transform -1 0 884 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_17
timestamp 1713260442
transform 1 0 884 0 1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_20
timestamp 1713260442
transform -1 0 940 0 1 505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_113
timestamp 1713260442
transform 1 0 940 0 1 505
box -2 -3 98 103
use FILL  FILL_5_1_0
timestamp 1713260442
transform -1 0 1044 0 1 505
box -2 -3 10 103
use FILL  FILL_5_1_1
timestamp 1713260442
transform -1 0 1052 0 1 505
box -2 -3 10 103
use OAI21X1  OAI21X1_68
timestamp 1713260442
transform -1 0 1084 0 1 505
box -2 -3 34 103
use INVX1  INVX1_14
timestamp 1713260442
transform -1 0 1100 0 1 505
box -2 -3 18 103
use NAND2X1  NAND2X1_36
timestamp 1713260442
transform 1 0 1100 0 1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_33
timestamp 1713260442
transform -1 0 1156 0 1 505
box -2 -3 34 103
use AOI21X1  AOI21X1_90
timestamp 1713260442
transform 1 0 1156 0 1 505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_89
timestamp 1713260442
transform -1 0 1284 0 1 505
box -2 -3 98 103
use OAI21X1  OAI21X1_156
timestamp 1713260442
transform 1 0 1284 0 1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_86
timestamp 1713260442
transform -1 0 1340 0 1 505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_63
timestamp 1713260442
transform 1 0 1340 0 1 505
box -2 -3 98 103
use BUFX4  BUFX4_27
timestamp 1713260442
transform 1 0 1436 0 1 505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_47
timestamp 1713260442
transform -1 0 1564 0 1 505
box -2 -3 98 103
use FILL  FILL_5_2_0
timestamp 1713260442
transform -1 0 1572 0 1 505
box -2 -3 10 103
use FILL  FILL_5_2_1
timestamp 1713260442
transform -1 0 1580 0 1 505
box -2 -3 10 103
use INVX1  INVX1_29
timestamp 1713260442
transform -1 0 1596 0 1 505
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_12
timestamp 1713260442
transform -1 0 1692 0 1 505
box -2 -3 98 103
use MUX2X1  MUX2X1_17
timestamp 1713260442
transform 1 0 1692 0 1 505
box -2 -3 50 103
use AOI21X1  AOI21X1_78
timestamp 1713260442
transform 1 0 1740 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_139
timestamp 1713260442
transform -1 0 1804 0 1 505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_52
timestamp 1713260442
transform 1 0 1804 0 1 505
box -2 -3 98 103
use INVX1  INVX1_27
timestamp 1713260442
transform 1 0 1900 0 1 505
box -2 -3 18 103
use NAND2X1  NAND2X1_79
timestamp 1713260442
transform -1 0 1940 0 1 505
box -2 -3 26 103
use AOI21X1  AOI21X1_99
timestamp 1713260442
transform 1 0 1940 0 1 505
box -2 -3 34 103
use NOR2X1  NOR2X1_74
timestamp 1713260442
transform -1 0 1996 0 1 505
box -2 -3 26 103
use NAND2X1  NAND2X1_73
timestamp 1713260442
transform -1 0 2020 0 1 505
box -2 -3 26 103
use AOI21X1  AOI21X1_98
timestamp 1713260442
transform -1 0 2052 0 1 505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_109
timestamp 1713260442
transform 1 0 4 0 -1 705
box -2 -3 98 103
use OAI21X1  OAI21X1_29
timestamp 1713260442
transform -1 0 132 0 -1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_32
timestamp 1713260442
transform -1 0 156 0 -1 705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_86
timestamp 1713260442
transform 1 0 156 0 -1 705
box -2 -3 98 103
use OAI21X1  OAI21X1_46
timestamp 1713260442
transform 1 0 252 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_150
timestamp 1713260442
transform 1 0 284 0 -1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_74
timestamp 1713260442
transform -1 0 340 0 -1 705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_57
timestamp 1713260442
transform 1 0 340 0 -1 705
box -2 -3 98 103
use OAI21X1  OAI21X1_147
timestamp 1713260442
transform 1 0 436 0 -1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_30
timestamp 1713260442
transform 1 0 468 0 -1 705
box -2 -3 34 103
use FILL  FILL_6_0_0
timestamp 1713260442
transform 1 0 500 0 -1 705
box -2 -3 10 103
use FILL  FILL_6_0_1
timestamp 1713260442
transform 1 0 508 0 -1 705
box -2 -3 10 103
use OAI21X1  OAI21X1_77
timestamp 1713260442
transform 1 0 516 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_65
timestamp 1713260442
transform -1 0 580 0 -1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_67
timestamp 1713260442
transform -1 0 604 0 -1 705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_20
timestamp 1713260442
transform 1 0 604 0 -1 705
box -2 -3 98 103
use AOI21X1  AOI21X1_87
timestamp 1713260442
transform 1 0 700 0 -1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_61
timestamp 1713260442
transform 1 0 732 0 -1 705
box -2 -3 26 103
use BUFX4  BUFX4_3
timestamp 1713260442
transform 1 0 756 0 -1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_68
timestamp 1713260442
transform -1 0 812 0 -1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_97
timestamp 1713260442
transform -1 0 844 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_111
timestamp 1713260442
transform -1 0 876 0 -1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_72
timestamp 1713260442
transform -1 0 900 0 -1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_141
timestamp 1713260442
transform -1 0 932 0 -1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_71
timestamp 1713260442
transform -1 0 956 0 -1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_130
timestamp 1713260442
transform -1 0 988 0 -1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_72
timestamp 1713260442
transform -1 0 1020 0 -1 705
box -2 -3 34 103
use FILL  FILL_6_1_0
timestamp 1713260442
transform -1 0 1028 0 -1 705
box -2 -3 10 103
use FILL  FILL_6_1_1
timestamp 1713260442
transform -1 0 1036 0 -1 705
box -2 -3 10 103
use OAI21X1  OAI21X1_133
timestamp 1713260442
transform -1 0 1068 0 -1 705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_80
timestamp 1713260442
transform 1 0 1068 0 -1 705
box -2 -3 98 103
use AOI21X1  AOI21X1_59
timestamp 1713260442
transform 1 0 1164 0 -1 705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_61
timestamp 1713260442
transform -1 0 1292 0 -1 705
box -2 -3 98 103
use AOI21X1  AOI21X1_9
timestamp 1713260442
transform -1 0 1324 0 -1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_82
timestamp 1713260442
transform 1 0 1324 0 -1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_154
timestamp 1713260442
transform -1 0 1380 0 -1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_73
timestamp 1713260442
transform 1 0 1380 0 -1 705
box -2 -3 34 103
use BUFX4  BUFX4_22
timestamp 1713260442
transform 1 0 1412 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_131
timestamp 1713260442
transform -1 0 1476 0 -1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_76
timestamp 1713260442
transform 1 0 1476 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_155
timestamp 1713260442
transform 1 0 1508 0 -1 705
box -2 -3 34 103
use FILL  FILL_6_2_0
timestamp 1713260442
transform 1 0 1540 0 -1 705
box -2 -3 10 103
use FILL  FILL_6_2_1
timestamp 1713260442
transform 1 0 1548 0 -1 705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_62
timestamp 1713260442
transform 1 0 1556 0 -1 705
box -2 -3 98 103
use MUX2X1  MUX2X1_20
timestamp 1713260442
transform 1 0 1652 0 -1 705
box -2 -3 50 103
use INVX1  INVX1_47
timestamp 1713260442
transform -1 0 1716 0 -1 705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_15
timestamp 1713260442
transform -1 0 1812 0 -1 705
box -2 -3 98 103
use MUX2X1  MUX2X1_3
timestamp 1713260442
transform -1 0 1860 0 -1 705
box -2 -3 50 103
use AOI21X1  AOI21X1_50
timestamp 1713260442
transform 1 0 1860 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_95
timestamp 1713260442
transform -1 0 1924 0 -1 705
box -2 -3 34 103
use INVX4  INVX4_4
timestamp 1713260442
transform 1 0 1924 0 -1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_128
timestamp 1713260442
transform -1 0 1980 0 -1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_70
timestamp 1713260442
transform 1 0 1980 0 -1 705
box -2 -3 26 103
use AOI21X1  AOI21X1_71
timestamp 1713260442
transform -1 0 2036 0 -1 705
box -2 -3 34 103
use FILL  FILL_7_1
timestamp 1713260442
transform -1 0 2044 0 -1 705
box -2 -3 10 103
use FILL  FILL_7_2
timestamp 1713260442
transform -1 0 2052 0 -1 705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_17
timestamp 1713260442
transform 1 0 4 0 1 705
box -2 -3 98 103
use NOR2X1  NOR2X1_59
timestamp 1713260442
transform 1 0 100 0 1 705
box -2 -3 26 103
use AOI21X1  AOI21X1_85
timestamp 1713260442
transform -1 0 156 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_22
timestamp 1713260442
transform -1 0 188 0 1 705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_118
timestamp 1713260442
transform 1 0 188 0 1 705
box -2 -3 98 103
use NAND2X1  NAND2X1_49
timestamp 1713260442
transform 1 0 284 0 1 705
box -2 -3 26 103
use INVX1  INVX1_56
timestamp 1713260442
transform -1 0 324 0 1 705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_111
timestamp 1713260442
transform 1 0 324 0 1 705
box -2 -3 98 103
use NAND2X1  NAND2X1_34
timestamp 1713260442
transform 1 0 420 0 1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_31
timestamp 1713260442
transform -1 0 476 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_114
timestamp 1713260442
transform 1 0 476 0 1 705
box -2 -3 34 103
use FILL  FILL_7_0_0
timestamp 1713260442
transform 1 0 508 0 1 705
box -2 -3 10 103
use FILL  FILL_7_0_1
timestamp 1713260442
transform 1 0 516 0 1 705
box -2 -3 10 103
use OAI21X1  OAI21X1_136
timestamp 1713260442
transform 1 0 524 0 1 705
box -2 -3 34 103
use BUFX4  BUFX4_6
timestamp 1713260442
transform -1 0 588 0 1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_52
timestamp 1713260442
transform -1 0 612 0 1 705
box -2 -3 26 103
use OAI22X1  OAI22X1_11
timestamp 1713260442
transform -1 0 652 0 1 705
box -2 -3 42 103
use OAI21X1  OAI21X1_138
timestamp 1713260442
transform 1 0 652 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_94
timestamp 1713260442
transform 1 0 684 0 1 705
box -2 -3 34 103
use OAI22X1  OAI22X1_7
timestamp 1713260442
transform -1 0 756 0 1 705
box -2 -3 42 103
use OAI22X1  OAI22X1_4
timestamp 1713260442
transform -1 0 796 0 1 705
box -2 -3 42 103
use OAI22X1  OAI22X1_13
timestamp 1713260442
transform -1 0 836 0 1 705
box -2 -3 42 103
use OAI21X1  OAI21X1_96
timestamp 1713260442
transform 1 0 836 0 1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_51
timestamp 1713260442
transform -1 0 900 0 1 705
box -2 -3 34 103
use OAI22X1  OAI22X1_12
timestamp 1713260442
transform 1 0 900 0 1 705
box -2 -3 42 103
use NOR2X1  NOR2X1_44
timestamp 1713260442
transform 1 0 940 0 1 705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_4
timestamp 1713260442
transform -1 0 1060 0 1 705
box -2 -3 98 103
use FILL  FILL_7_1_0
timestamp 1713260442
transform 1 0 1060 0 1 705
box -2 -3 10 103
use FILL  FILL_7_1_1
timestamp 1713260442
transform 1 0 1068 0 1 705
box -2 -3 10 103
use NAND2X1  NAND2X1_93
timestamp 1713260442
transform 1 0 1076 0 1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_161
timestamp 1713260442
transform -1 0 1132 0 1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_54
timestamp 1713260442
transform 1 0 1132 0 1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_148
timestamp 1713260442
transform -1 0 1188 0 1 705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_32
timestamp 1713260442
transform -1 0 1284 0 1 705
box -2 -3 98 103
use NOR2X1  NOR2X1_11
timestamp 1713260442
transform 1 0 1284 0 1 705
box -2 -3 26 103
use NOR2X1  NOR2X1_25
timestamp 1713260442
transform 1 0 1308 0 1 705
box -2 -3 26 103
use AOI21X1  AOI21X1_21
timestamp 1713260442
transform -1 0 1364 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_15
timestamp 1713260442
transform 1 0 1364 0 1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_18
timestamp 1713260442
transform -1 0 1420 0 1 705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_127
timestamp 1713260442
transform 1 0 1420 0 1 705
box -2 -3 98 103
use FILL  FILL_7_2_0
timestamp 1713260442
transform 1 0 1516 0 1 705
box -2 -3 10 103
use FILL  FILL_7_2_1
timestamp 1713260442
transform 1 0 1524 0 1 705
box -2 -3 10 103
use AOI21X1  AOI21X1_77
timestamp 1713260442
transform 1 0 1532 0 1 705
box -2 -3 34 103
use INVX1  INVX1_50
timestamp 1713260442
transform 1 0 1564 0 1 705
box -2 -3 18 103
use OAI21X1  OAI21X1_135
timestamp 1713260442
transform -1 0 1612 0 1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_84
timestamp 1713260442
transform -1 0 1636 0 1 705
box -2 -3 26 103
use NOR2X1  NOR2X1_19
timestamp 1713260442
transform 1 0 1636 0 1 705
box -2 -3 26 103
use AOI21X1  AOI21X1_16
timestamp 1713260442
transform -1 0 1692 0 1 705
box -2 -3 34 103
use BUFX4  BUFX4_31
timestamp 1713260442
transform 1 0 1692 0 1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_54
timestamp 1713260442
transform -1 0 1756 0 1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_7
timestamp 1713260442
transform 1 0 1756 0 1 705
box -2 -3 26 103
use AOI21X1  AOI21X1_5
timestamp 1713260442
transform -1 0 1812 0 1 705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_76
timestamp 1713260442
transform -1 0 1908 0 1 705
box -2 -3 98 103
use INVX1  INVX1_15
timestamp 1713260442
transform -1 0 1924 0 1 705
box -2 -3 18 103
use AOI21X1  AOI21X1_95
timestamp 1713260442
transform 1 0 1924 0 1 705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_68
timestamp 1713260442
transform -1 0 2052 0 1 705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_112
timestamp 1713260442
transform -1 0 100 0 -1 905
box -2 -3 98 103
use NAND2X1  NAND2X1_35
timestamp 1713260442
transform 1 0 100 0 -1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_32
timestamp 1713260442
transform -1 0 156 0 -1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_25
timestamp 1713260442
transform -1 0 180 0 -1 905
box -2 -3 26 103
use AOI21X1  AOI21X1_83
timestamp 1713260442
transform 1 0 180 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_146
timestamp 1713260442
transform -1 0 244 0 -1 905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_44
timestamp 1713260442
transform 1 0 244 0 -1 905
box -2 -3 98 103
use NOR2X1  NOR2X1_16
timestamp 1713260442
transform 1 0 340 0 -1 905
box -2 -3 26 103
use AOI21X1  AOI21X1_13
timestamp 1713260442
transform -1 0 396 0 -1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_55
timestamp 1713260442
transform 1 0 396 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_102
timestamp 1713260442
transform -1 0 460 0 -1 905
box -2 -3 34 103
use INVX1  INVX1_32
timestamp 1713260442
transform -1 0 476 0 -1 905
box -2 -3 18 103
use FILL  FILL_8_0_0
timestamp 1713260442
transform -1 0 484 0 -1 905
box -2 -3 10 103
use FILL  FILL_8_0_1
timestamp 1713260442
transform -1 0 492 0 -1 905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_124
timestamp 1713260442
transform -1 0 588 0 -1 905
box -2 -3 98 103
use NAND2X1  NAND2X1_15
timestamp 1713260442
transform 1 0 588 0 -1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_12
timestamp 1713260442
transform -1 0 644 0 -1 905
box -2 -3 34 103
use BUFX4  BUFX4_30
timestamp 1713260442
transform 1 0 644 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_116
timestamp 1713260442
transform -1 0 708 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_137
timestamp 1713260442
transform -1 0 740 0 -1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_56
timestamp 1713260442
transform -1 0 772 0 -1 905
box -2 -3 34 103
use BUFX4  BUFX4_19
timestamp 1713260442
transform -1 0 804 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_104
timestamp 1713260442
transform 1 0 804 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_73
timestamp 1713260442
transform -1 0 868 0 -1 905
box -2 -3 34 103
use INVX8  INVX8_3
timestamp 1713260442
transform 1 0 868 0 -1 905
box -2 -3 42 103
use AOI21X1  AOI21X1_79
timestamp 1713260442
transform 1 0 908 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_129
timestamp 1713260442
transform -1 0 972 0 -1 905
box -2 -3 34 103
use INVX1  INVX1_46
timestamp 1713260442
transform -1 0 988 0 -1 905
box -2 -3 18 103
use NAND2X1  NAND2X1_97
timestamp 1713260442
transform 1 0 988 0 -1 905
box -2 -3 26 103
use FILL  FILL_8_1_0
timestamp 1713260442
transform -1 0 1020 0 -1 905
box -2 -3 10 103
use FILL  FILL_8_1_1
timestamp 1713260442
transform -1 0 1028 0 -1 905
box -2 -3 10 103
use OAI21X1  OAI21X1_165
timestamp 1713260442
transform -1 0 1060 0 -1 905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_8
timestamp 1713260442
transform -1 0 1156 0 -1 905
box -2 -3 98 103
use AOI21X1  AOI21X1_75
timestamp 1713260442
transform -1 0 1188 0 -1 905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_79
timestamp 1713260442
transform -1 0 1284 0 -1 905
box -2 -3 98 103
use NOR2X1  NOR2X1_10
timestamp 1713260442
transform 1 0 1284 0 -1 905
box -2 -3 26 103
use AOI21X1  AOI21X1_8
timestamp 1713260442
transform -1 0 1340 0 -1 905
box -2 -3 34 103
use BUFX4  BUFX4_1
timestamp 1713260442
transform 1 0 1340 0 -1 905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_106
timestamp 1713260442
transform -1 0 1468 0 -1 905
box -2 -3 98 103
use OAI21X1  OAI21X1_134
timestamp 1713260442
transform -1 0 1500 0 -1 905
box -2 -3 34 103
use MUX2X1  MUX2X1_11
timestamp 1713260442
transform 1 0 1500 0 -1 905
box -2 -3 50 103
use FILL  FILL_8_2_0
timestamp 1713260442
transform -1 0 1556 0 -1 905
box -2 -3 10 103
use FILL  FILL_8_2_1
timestamp 1713260442
transform -1 0 1564 0 -1 905
box -2 -3 10 103
use AOI21X1  AOI21X1_38
timestamp 1713260442
transform -1 0 1596 0 -1 905
box -2 -3 34 103
use INVX1  INVX1_49
timestamp 1713260442
transform -1 0 1612 0 -1 905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_31
timestamp 1713260442
transform -1 0 1708 0 -1 905
box -2 -3 98 103
use OAI21X1  OAI21X1_101
timestamp 1713260442
transform 1 0 1708 0 -1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_28
timestamp 1713260442
transform -1 0 1764 0 -1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_25
timestamp 1713260442
transform -1 0 1796 0 -1 905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_105
timestamp 1713260442
transform -1 0 1892 0 -1 905
box -2 -3 98 103
use MUX2X1  MUX2X1_6
timestamp 1713260442
transform -1 0 1940 0 -1 905
box -2 -3 50 103
use INVX1  INVX1_45
timestamp 1713260442
transform -1 0 1956 0 -1 905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_55
timestamp 1713260442
transform -1 0 2052 0 -1 905
box -2 -3 98 103
use CLKBUF1  CLKBUF1_4
timestamp 1713260442
transform 1 0 4 0 1 905
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_1
timestamp 1713260442
transform 1 0 76 0 1 905
box -2 -3 98 103
use OAI21X1  OAI21X1_158
timestamp 1713260442
transform 1 0 172 0 1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_90
timestamp 1713260442
transform 1 0 204 0 1 905
box -2 -3 26 103
use AOI21X1  AOI21X1_68
timestamp 1713260442
transform 1 0 228 0 1 905
box -2 -3 34 103
use INVX1  INVX1_44
timestamp 1713260442
transform 1 0 260 0 1 905
box -2 -3 18 103
use AOI21X1  AOI21X1_84
timestamp 1713260442
transform 1 0 276 0 1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_29
timestamp 1713260442
transform 1 0 308 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_63
timestamp 1713260442
transform 1 0 340 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_66
timestamp 1713260442
transform 1 0 372 0 1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_31
timestamp 1713260442
transform -1 0 436 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_67
timestamp 1713260442
transform -1 0 468 0 1 905
box -2 -3 34 103
use OAI22X1  OAI22X1_14
timestamp 1713260442
transform 1 0 468 0 1 905
box -2 -3 42 103
use FILL  FILL_9_0_0
timestamp 1713260442
transform -1 0 516 0 1 905
box -2 -3 10 103
use FILL  FILL_9_0_1
timestamp 1713260442
transform -1 0 524 0 1 905
box -2 -3 10 103
use BUFX4  BUFX4_20
timestamp 1713260442
transform -1 0 556 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_64
timestamp 1713260442
transform -1 0 588 0 1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_32
timestamp 1713260442
transform 1 0 588 0 1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_39
timestamp 1713260442
transform -1 0 652 0 1 905
box -2 -3 34 103
use BUFX4  BUFX4_21
timestamp 1713260442
transform 1 0 652 0 1 905
box -2 -3 34 103
use INVX8  INVX8_4
timestamp 1713260442
transform -1 0 724 0 1 905
box -2 -3 42 103
use OAI22X1  OAI22X1_6
timestamp 1713260442
transform -1 0 764 0 1 905
box -2 -3 42 103
use OAI21X1  OAI21X1_82
timestamp 1713260442
transform -1 0 796 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_149
timestamp 1713260442
transform -1 0 828 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_105
timestamp 1713260442
transform -1 0 860 0 1 905
box -2 -3 34 103
use OAI22X1  OAI22X1_5
timestamp 1713260442
transform 1 0 860 0 1 905
box -2 -3 42 103
use AOI21X1  AOI21X1_58
timestamp 1713260442
transform -1 0 932 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_140
timestamp 1713260442
transform -1 0 964 0 1 905
box -2 -3 34 103
use BUFX4  BUFX4_18
timestamp 1713260442
transform -1 0 996 0 1 905
box -2 -3 34 103
use BUFX4  BUFX4_43
timestamp 1713260442
transform -1 0 1028 0 1 905
box -2 -3 34 103
use FILL  FILL_9_1_0
timestamp 1713260442
transform 1 0 1028 0 1 905
box -2 -3 10 103
use FILL  FILL_9_1_1
timestamp 1713260442
transform 1 0 1036 0 1 905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_108
timestamp 1713260442
transform 1 0 1044 0 1 905
box -2 -3 98 103
use OAI21X1  OAI21X1_103
timestamp 1713260442
transform 1 0 1140 0 1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_31
timestamp 1713260442
transform 1 0 1172 0 1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_28
timestamp 1713260442
transform -1 0 1228 0 1 905
box -2 -3 34 103
use BUFX4  BUFX4_2
timestamp 1713260442
transform -1 0 1260 0 1 905
box -2 -3 34 103
use BUFX4  BUFX4_39
timestamp 1713260442
transform 1 0 1260 0 1 905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_41
timestamp 1713260442
transform 1 0 1292 0 1 905
box -2 -3 98 103
use AOI21X1  AOI21X1_10
timestamp 1713260442
transform 1 0 1388 0 1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_13
timestamp 1713260442
transform -1 0 1444 0 1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_71
timestamp 1713260442
transform 1 0 1444 0 1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_37
timestamp 1713260442
transform 1 0 1476 0 1 905
box -2 -3 34 103
use BUFX4  BUFX4_23
timestamp 1713260442
transform 1 0 1508 0 1 905
box -2 -3 34 103
use FILL  FILL_9_2_0
timestamp 1713260442
transform -1 0 1548 0 1 905
box -2 -3 10 103
use FILL  FILL_9_2_1
timestamp 1713260442
transform -1 0 1556 0 1 905
box -2 -3 10 103
use OR2X2  OR2X2_1
timestamp 1713260442
transform -1 0 1588 0 1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_35
timestamp 1713260442
transform -1 0 1620 0 1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_29
timestamp 1713260442
transform 1 0 1620 0 1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_26
timestamp 1713260442
transform -1 0 1676 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_109
timestamp 1713260442
transform -1 0 1708 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_69
timestamp 1713260442
transform 1 0 1708 0 1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_34
timestamp 1713260442
transform -1 0 1772 0 1 905
box -2 -3 34 103
use MUX2X1  MUX2X1_9
timestamp 1713260442
transform 1 0 1772 0 1 905
box -2 -3 50 103
use INVX1  INVX1_35
timestamp 1713260442
transform -1 0 1836 0 1 905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_13
timestamp 1713260442
transform -1 0 1932 0 1 905
box -2 -3 98 103
use INVX1  INVX1_31
timestamp 1713260442
transform -1 0 1948 0 1 905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_28
timestamp 1713260442
transform -1 0 2044 0 1 905
box -2 -3 98 103
use FILL  FILL_10_1
timestamp 1713260442
transform 1 0 2044 0 1 905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_94
timestamp 1713260442
transform -1 0 100 0 -1 1105
box -2 -3 98 103
use INVX1  INVX1_13
timestamp 1713260442
transform 1 0 100 0 -1 1105
box -2 -3 18 103
use OAI21X1  OAI21X1_38
timestamp 1713260442
transform 1 0 116 0 -1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_41
timestamp 1713260442
transform -1 0 172 0 -1 1105
box -2 -3 26 103
use MUX2X1  MUX2X1_22
timestamp 1713260442
transform -1 0 220 0 -1 1105
box -2 -3 50 103
use INVX1  INVX1_43
timestamp 1713260442
transform 1 0 220 0 -1 1105
box -2 -3 18 103
use OAI21X1  OAI21X1_123
timestamp 1713260442
transform 1 0 236 0 -1 1105
box -2 -3 34 103
use INVX1  INVX1_55
timestamp 1713260442
transform 1 0 268 0 -1 1105
box -2 -3 18 103
use AOI21X1  AOI21X1_69
timestamp 1713260442
transform 1 0 284 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_124
timestamp 1713260442
transform -1 0 348 0 -1 1105
box -2 -3 34 103
use INVX1  INVX1_11
timestamp 1713260442
transform 1 0 348 0 -1 1105
box -2 -3 18 103
use OAI21X1  OAI21X1_145
timestamp 1713260442
transform 1 0 364 0 -1 1105
box -2 -3 34 103
use AOI21X1  AOI21X1_82
timestamp 1713260442
transform -1 0 428 0 -1 1105
box -2 -3 34 103
use AOI21X1  AOI21X1_70
timestamp 1713260442
transform 1 0 428 0 -1 1105
box -2 -3 34 103
use BUFX4  BUFX4_5
timestamp 1713260442
transform -1 0 492 0 -1 1105
box -2 -3 34 103
use FILL  FILL_10_0_0
timestamp 1713260442
transform 1 0 492 0 -1 1105
box -2 -3 10 103
use FILL  FILL_10_0_1
timestamp 1713260442
transform 1 0 500 0 -1 1105
box -2 -3 10 103
use BUFX4  BUFX4_4
timestamp 1713260442
transform 1 0 508 0 -1 1105
box -2 -3 34 103
use BUFX4  BUFX4_32
timestamp 1713260442
transform -1 0 572 0 -1 1105
box -2 -3 34 103
use OAI22X1  OAI22X1_2
timestamp 1713260442
transform -1 0 612 0 -1 1105
box -2 -3 42 103
use BUFX4  BUFX4_37
timestamp 1713260442
transform -1 0 644 0 -1 1105
box -2 -3 34 103
use INVX1  INVX1_28
timestamp 1713260442
transform 1 0 644 0 -1 1105
box -2 -3 18 103
use AOI21X1  AOI21X1_45
timestamp 1713260442
transform -1 0 692 0 -1 1105
box -2 -3 34 103
use OAI22X1  OAI22X1_8
timestamp 1713260442
transform 1 0 692 0 -1 1105
box -2 -3 42 103
use NOR2X1  NOR2X1_49
timestamp 1713260442
transform 1 0 732 0 -1 1105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_116
timestamp 1713260442
transform 1 0 756 0 -1 1105
box -2 -3 98 103
use NAND2X1  NAND2X1_69
timestamp 1713260442
transform -1 0 876 0 -1 1105
box -2 -3 26 103
use NOR2X1  NOR2X1_46
timestamp 1713260442
transform -1 0 900 0 -1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_108
timestamp 1713260442
transform -1 0 932 0 -1 1105
box -2 -3 34 103
use BUFX4  BUFX4_40
timestamp 1713260442
transform -1 0 964 0 -1 1105
box -2 -3 34 103
use INVX1  INVX1_52
timestamp 1713260442
transform -1 0 980 0 -1 1105
box -2 -3 18 103
use NAND2X1  NAND2X1_7
timestamp 1713260442
transform 1 0 980 0 -1 1105
box -2 -3 26 103
use FILL  FILL_10_1_0
timestamp 1713260442
transform -1 0 1012 0 -1 1105
box -2 -3 10 103
use FILL  FILL_10_1_1
timestamp 1713260442
transform -1 0 1020 0 -1 1105
box -2 -3 10 103
use OAI21X1  OAI21X1_7
timestamp 1713260442
transform -1 0 1052 0 -1 1105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_39
timestamp 1713260442
transform -1 0 1148 0 -1 1105
box -2 -3 98 103
use BUFX4  BUFX4_16
timestamp 1713260442
transform 1 0 1148 0 -1 1105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_77
timestamp 1713260442
transform 1 0 1180 0 -1 1105
box -2 -3 98 103
use NOR2X1  NOR2X1_8
timestamp 1713260442
transform 1 0 1276 0 -1 1105
box -2 -3 26 103
use AOI21X1  AOI21X1_6
timestamp 1713260442
transform -1 0 1332 0 -1 1105
box -2 -3 34 103
use MUX2X1  MUX2X1_10
timestamp 1713260442
transform 1 0 1332 0 -1 1105
box -2 -3 50 103
use INVX1  INVX1_37
timestamp 1713260442
transform -1 0 1396 0 -1 1105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_29
timestamp 1713260442
transform -1 0 1492 0 -1 1105
box -2 -3 98 103
use FILL  FILL_10_2_0
timestamp 1713260442
transform 1 0 1492 0 -1 1105
box -2 -3 10 103
use FILL  FILL_10_2_1
timestamp 1713260442
transform 1 0 1500 0 -1 1105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_69
timestamp 1713260442
transform 1 0 1508 0 -1 1105
box -2 -3 98 103
use AOI21X1  AOI21X1_96
timestamp 1713260442
transform 1 0 1604 0 -1 1105
box -2 -3 34 103
use NOR2X1  NOR2X1_71
timestamp 1713260442
transform -1 0 1660 0 -1 1105
box -2 -3 26 103
use AOI21X1  AOI21X1_57
timestamp 1713260442
transform 1 0 1660 0 -1 1105
box -2 -3 34 103
use BUFX4  BUFX4_28
timestamp 1713260442
transform 1 0 1692 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_106
timestamp 1713260442
transform -1 0 1756 0 -1 1105
box -2 -3 34 103
use INVX1  INVX1_33
timestamp 1713260442
transform -1 0 1772 0 -1 1105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_53
timestamp 1713260442
transform -1 0 1868 0 -1 1105
box -2 -3 98 103
use MUX2X1  MUX2X1_18
timestamp 1713260442
transform 1 0 1868 0 -1 1105
box -2 -3 50 103
use MUX2X1  MUX2X1_4
timestamp 1713260442
transform 1 0 1916 0 -1 1105
box -2 -3 50 103
use OAI21X1  OAI21X1_41
timestamp 1713260442
transform 1 0 1964 0 -1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_44
timestamp 1713260442
transform -1 0 2020 0 -1 1105
box -2 -3 26 103
use NAND2X1  NAND2X1_81
timestamp 1713260442
transform -1 0 2044 0 -1 1105
box -2 -3 26 103
use FILL  FILL_11_1
timestamp 1713260442
transform -1 0 2052 0 -1 1105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_97
timestamp 1713260442
transform 1 0 4 0 1 1105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_98
timestamp 1713260442
transform 1 0 100 0 1 1105
box -2 -3 98 103
use INVX1  INVX1_21
timestamp 1713260442
transform 1 0 196 0 1 1105
box -2 -3 18 103
use MUX2X1  MUX2X1_23
timestamp 1713260442
transform 1 0 212 0 1 1105
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_33
timestamp 1713260442
transform 1 0 260 0 1 1105
box -2 -3 98 103
use NAND2X1  NAND2X1_1
timestamp 1713260442
transform 1 0 356 0 1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_1
timestamp 1713260442
transform -1 0 412 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_76
timestamp 1713260442
transform 1 0 412 0 1 1105
box -2 -3 34 103
use AOI21X1  AOI21X1_43
timestamp 1713260442
transform -1 0 476 0 1 1105
box -2 -3 34 103
use BUFX4  BUFX4_44
timestamp 1713260442
transform -1 0 508 0 1 1105
box -2 -3 34 103
use FILL  FILL_11_0_0
timestamp 1713260442
transform 1 0 508 0 1 1105
box -2 -3 10 103
use FILL  FILL_11_0_1
timestamp 1713260442
transform 1 0 516 0 1 1105
box -2 -3 10 103
use OAI21X1  OAI21X1_4
timestamp 1713260442
transform 1 0 524 0 1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_4
timestamp 1713260442
transform -1 0 580 0 1 1105
box -2 -3 26 103
use AOI21X1  AOI21X1_46
timestamp 1713260442
transform -1 0 612 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_79
timestamp 1713260442
transform 1 0 612 0 1 1105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_36
timestamp 1713260442
transform -1 0 740 0 1 1105
box -2 -3 98 103
use BUFX4  BUFX4_36
timestamp 1713260442
transform -1 0 772 0 1 1105
box -2 -3 34 103
use BUFX4  BUFX4_35
timestamp 1713260442
transform 1 0 772 0 1 1105
box -2 -3 34 103
use BUFX4  BUFX4_34
timestamp 1713260442
transform 1 0 804 0 1 1105
box -2 -3 34 103
use AOI21X1  AOI21X1_63
timestamp 1713260442
transform -1 0 868 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_20
timestamp 1713260442
transform 1 0 868 0 1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_23
timestamp 1713260442
transform 1 0 900 0 1 1105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_40
timestamp 1713260442
transform 1 0 924 0 1 1105
box -2 -3 98 103
use FILL  FILL_11_1_0
timestamp 1713260442
transform 1 0 1020 0 1 1105
box -2 -3 10 103
use FILL  FILL_11_1_1
timestamp 1713260442
transform 1 0 1028 0 1 1105
box -2 -3 10 103
use NAND2X1  NAND2X1_8
timestamp 1713260442
transform 1 0 1036 0 1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_8
timestamp 1713260442
transform -1 0 1092 0 1 1105
box -2 -3 34 103
use BUFX4  BUFX4_47
timestamp 1713260442
transform 1 0 1092 0 1 1105
box -2 -3 34 103
use XNOR2X1  XNOR2X1_2
timestamp 1713260442
transform -1 0 1180 0 1 1105
box -2 -3 58 103
use BUFX4  BUFX4_17
timestamp 1713260442
transform -1 0 1212 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_126
timestamp 1713260442
transform -1 0 1244 0 1 1105
box -2 -3 34 103
use AOI21X1  AOI21X1_61
timestamp 1713260442
transform 1 0 1244 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_112
timestamp 1713260442
transform -1 0 1308 0 1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_56
timestamp 1713260442
transform 1 0 1308 0 1 1105
box -2 -3 26 103
use DFFSR  DFFSR_2
timestamp 1713260442
transform -1 0 1508 0 1 1105
box -2 -3 178 103
use NOR2X1  NOR2X1_31
timestamp 1713260442
transform -1 0 1532 0 1 1105
box -2 -3 26 103
use FILL  FILL_11_2_0
timestamp 1713260442
transform -1 0 1540 0 1 1105
box -2 -3 10 103
use FILL  FILL_11_2_1
timestamp 1713260442
transform -1 0 1548 0 1 1105
box -2 -3 10 103
use AOI21X1  AOI21X1_22
timestamp 1713260442
transform -1 0 1580 0 1 1105
box -2 -3 34 103
use AOI21X1  AOI21X1_23
timestamp 1713260442
transform -1 0 1612 0 1 1105
box -2 -3 34 103
use NAND3X1  NAND3X1_8
timestamp 1713260442
transform -1 0 1644 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_51
timestamp 1713260442
transform 1 0 1644 0 1 1105
box -2 -3 34 103
use DFFSR  DFFSR_3
timestamp 1713260442
transform 1 0 1676 0 1 1105
box -2 -3 178 103
use DFFPOSX1  DFFPOSX1_81
timestamp 1713260442
transform -1 0 1948 0 1 1105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_54
timestamp 1713260442
transform 1 0 1948 0 1 1105
box -2 -3 98 103
use FILL  FILL_12_1
timestamp 1713260442
transform 1 0 2044 0 1 1105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_102
timestamp 1713260442
transform 1 0 4 0 -1 1305
box -2 -3 98 103
use INVX1  INVX1_42
timestamp 1713260442
transform 1 0 100 0 -1 1305
box -2 -3 18 103
use MUX2X1  MUX2X1_27
timestamp 1713260442
transform -1 0 164 0 -1 1305
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_114
timestamp 1713260442
transform 1 0 164 0 -1 1305
box -2 -3 98 103
use OAI21X1  OAI21X1_18
timestamp 1713260442
transform 1 0 260 0 -1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_21
timestamp 1713260442
transform -1 0 316 0 -1 1305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_120
timestamp 1713260442
transform 1 0 316 0 -1 1305
box -2 -3 98 103
use NAND2X1  NAND2X1_27
timestamp 1713260442
transform 1 0 412 0 -1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_121
timestamp 1713260442
transform 1 0 436 0 -1 1305
box -2 -3 34 103
use OAI22X1  OAI22X1_10
timestamp 1713260442
transform 1 0 468 0 -1 1305
box -2 -3 42 103
use FILL  FILL_12_0_0
timestamp 1713260442
transform 1 0 508 0 -1 1305
box -2 -3 10 103
use FILL  FILL_12_0_1
timestamp 1713260442
transform 1 0 516 0 -1 1305
box -2 -3 10 103
use AOI21X1  AOI21X1_44
timestamp 1713260442
transform 1 0 524 0 -1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_122
timestamp 1713260442
transform -1 0 588 0 -1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_70
timestamp 1713260442
transform -1 0 612 0 -1 1305
box -2 -3 26 103
use INVX1  INVX1_23
timestamp 1713260442
transform 1 0 612 0 -1 1305
box -2 -3 18 103
use OAI21X1  OAI21X1_78
timestamp 1713260442
transform -1 0 660 0 -1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_119
timestamp 1713260442
transform 1 0 660 0 -1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_45
timestamp 1713260442
transform 1 0 692 0 -1 1305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_85
timestamp 1713260442
transform -1 0 820 0 -1 1305
box -2 -3 98 103
use OAI21X1  OAI21X1_113
timestamp 1713260442
transform -1 0 852 0 -1 1305
box -2 -3 34 103
use NOR2X1  NOR2X1_47
timestamp 1713260442
transform -1 0 876 0 -1 1305
box -2 -3 26 103
use INVX1  INVX1_38
timestamp 1713260442
transform -1 0 892 0 -1 1305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_125
timestamp 1713260442
transform -1 0 988 0 -1 1305
box -2 -3 98 103
use NAND2X1  NAND2X1_16
timestamp 1713260442
transform 1 0 988 0 -1 1305
box -2 -3 26 103
use FILL  FILL_12_1_0
timestamp 1713260442
transform -1 0 1020 0 -1 1305
box -2 -3 10 103
use FILL  FILL_12_1_1
timestamp 1713260442
transform -1 0 1028 0 -1 1305
box -2 -3 10 103
use OAI21X1  OAI21X1_13
timestamp 1713260442
transform -1 0 1060 0 -1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_127
timestamp 1713260442
transform -1 0 1092 0 -1 1305
box -2 -3 34 103
use OAI22X1  OAI22X1_9
timestamp 1713260442
transform -1 0 1132 0 -1 1305
box -2 -3 42 103
use NOR2X1  NOR2X1_51
timestamp 1713260442
transform -1 0 1156 0 -1 1305
box -2 -3 26 103
use NOR2X1  NOR2X1_50
timestamp 1713260442
transform 1 0 1156 0 -1 1305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_126
timestamp 1713260442
transform -1 0 1276 0 -1 1305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_121
timestamp 1713260442
transform 1 0 1276 0 -1 1305
box -2 -3 98 103
use OAI21X1  OAI21X1_9
timestamp 1713260442
transform 1 0 1372 0 -1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_12
timestamp 1713260442
transform -1 0 1428 0 -1 1305
box -2 -3 26 103
use INVX1  INVX1_17
timestamp 1713260442
transform 1 0 1428 0 -1 1305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_30
timestamp 1713260442
transform -1 0 1540 0 -1 1305
box -2 -3 98 103
use FILL  FILL_12_2_0
timestamp 1713260442
transform 1 0 1540 0 -1 1305
box -2 -3 10 103
use FILL  FILL_12_2_1
timestamp 1713260442
transform 1 0 1548 0 -1 1305
box -2 -3 10 103
use NOR2X1  NOR2X1_24
timestamp 1713260442
transform 1 0 1556 0 -1 1305
box -2 -3 26 103
use AOI21X1  AOI21X1_20
timestamp 1713260442
transform -1 0 1612 0 -1 1305
box -2 -3 34 103
use AOI21X1  AOI21X1_66
timestamp 1713260442
transform -1 0 1644 0 -1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_120
timestamp 1713260442
transform -1 0 1676 0 -1 1305
box -2 -3 34 103
use AOI21X1  AOI21X1_64
timestamp 1713260442
transform 1 0 1676 0 -1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_117
timestamp 1713260442
transform -1 0 1740 0 -1 1305
box -2 -3 34 103
use BUFX4  BUFX4_10
timestamp 1713260442
transform 1 0 1740 0 -1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_83
timestamp 1713260442
transform -1 0 1796 0 -1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_85
timestamp 1713260442
transform -1 0 1820 0 -1 1305
box -2 -3 26 103
use BUFX4  BUFX4_8
timestamp 1713260442
transform 1 0 1820 0 -1 1305
box -2 -3 34 103
use INVX4  INVX4_6
timestamp 1713260442
transform 1 0 1852 0 -1 1305
box -2 -3 26 103
use INVX4  INVX4_8
timestamp 1713260442
transform -1 0 1900 0 -1 1305
box -2 -3 26 103
use INVX4  INVX4_7
timestamp 1713260442
transform 1 0 1900 0 -1 1305
box -2 -3 26 103
use MUX2X1  MUX2X1_5
timestamp 1713260442
transform 1 0 1924 0 -1 1305
box -2 -3 50 103
use AOI21X1  AOI21X1_97
timestamp 1713260442
transform 1 0 1972 0 -1 1305
box -2 -3 34 103
use INVX1  INVX1_39
timestamp 1713260442
transform -1 0 2020 0 -1 1305
box -2 -3 18 103
use NOR2X1  NOR2X1_72
timestamp 1713260442
transform 1 0 2020 0 -1 1305
box -2 -3 26 103
use FILL  FILL_13_1
timestamp 1713260442
transform -1 0 2052 0 -1 1305
box -2 -3 10 103
use DFFSR  DFFSR_10
timestamp 1713260442
transform -1 0 180 0 1 1305
box -2 -3 178 103
use NAND2X1  NAND2X1_33
timestamp 1713260442
transform -1 0 204 0 1 1305
box -2 -3 26 103
use DFFSR  DFFSR_16
timestamp 1713260442
transform -1 0 380 0 1 1305
box -2 -3 178 103
use OAI21X1  OAI21X1_24
timestamp 1713260442
transform 1 0 380 0 1 1305
box -2 -3 34 103
use AOI21X1  AOI21X1_67
timestamp 1713260442
transform 1 0 412 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_118
timestamp 1713260442
transform -1 0 476 0 1 1305
box -2 -3 34 103
use AOI21X1  AOI21X1_65
timestamp 1713260442
transform -1 0 508 0 1 1305
box -2 -3 34 103
use FILL  FILL_13_0_0
timestamp 1713260442
transform 1 0 508 0 1 1305
box -2 -3 10 103
use FILL  FILL_13_0_1
timestamp 1713260442
transform 1 0 516 0 1 1305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_82
timestamp 1713260442
transform 1 0 524 0 1 1305
box -2 -3 98 103
use NAND2X1  NAND2X1_45
timestamp 1713260442
transform 1 0 620 0 1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_42
timestamp 1713260442
transform -1 0 676 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_125
timestamp 1713260442
transform 1 0 676 0 1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_48
timestamp 1713260442
transform -1 0 732 0 1 1305
box -2 -3 26 103
use AOI21X1  AOI21X1_62
timestamp 1713260442
transform 1 0 732 0 1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_57
timestamp 1713260442
transform 1 0 764 0 1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_52
timestamp 1713260442
transform -1 0 820 0 1 1305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_84
timestamp 1713260442
transform -1 0 916 0 1 1305
box -2 -3 98 103
use NAND2X1  NAND2X1_47
timestamp 1713260442
transform 1 0 916 0 1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_44
timestamp 1713260442
transform -1 0 972 0 1 1305
box -2 -3 34 103
use BUFX4  BUFX4_41
timestamp 1713260442
transform -1 0 1004 0 1 1305
box -2 -3 34 103
use FILL  FILL_13_1_0
timestamp 1713260442
transform 1 0 1004 0 1 1305
box -2 -3 10 103
use FILL  FILL_13_1_1
timestamp 1713260442
transform 1 0 1012 0 1 1305
box -2 -3 10 103
use BUFX4  BUFX4_42
timestamp 1713260442
transform 1 0 1020 0 1 1305
box -2 -3 34 103
use MUX2X1  MUX2X1_12
timestamp 1713260442
transform 1 0 1052 0 1 1305
box -2 -3 50 103
use OAI21X1  OAI21X1_14
timestamp 1713260442
transform 1 0 1100 0 1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_17
timestamp 1713260442
transform -1 0 1156 0 1 1305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_78
timestamp 1713260442
transform -1 0 1252 0 1 1305
box -2 -3 98 103
use NAND2X1  NAND2X1_98
timestamp 1713260442
transform -1 0 1276 0 1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_9
timestamp 1713260442
transform 1 0 1276 0 1 1305
box -2 -3 26 103
use NOR2X1  NOR2X1_3
timestamp 1713260442
transform 1 0 1300 0 1 1305
box -2 -3 26 103
use NOR2X1  NOR2X1_75
timestamp 1713260442
transform 1 0 1324 0 1 1305
box -2 -3 26 103
use NOR2X1  NOR2X1_9
timestamp 1713260442
transform 1 0 1348 0 1 1305
box -2 -3 26 103
use AOI21X1  AOI21X1_7
timestamp 1713260442
transform -1 0 1404 0 1 1305
box -2 -3 34 103
use BUFX4  BUFX4_9
timestamp 1713260442
transform -1 0 1436 0 1 1305
box -2 -3 34 103
use BUFX4  BUFX4_38
timestamp 1713260442
transform 1 0 1436 0 1 1305
box -2 -3 34 103
use BUFX4  BUFX4_7
timestamp 1713260442
transform 1 0 1468 0 1 1305
box -2 -3 34 103
use FILL  FILL_13_2_0
timestamp 1713260442
transform 1 0 1500 0 1 1305
box -2 -3 10 103
use FILL  FILL_13_2_1
timestamp 1713260442
transform 1 0 1508 0 1 1305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_14
timestamp 1713260442
transform 1 0 1516 0 1 1305
box -2 -3 98 103
use NOR2X1  NOR2X1_30
timestamp 1713260442
transform -1 0 1636 0 1 1305
box -2 -3 26 103
use INVX1  INVX1_41
timestamp 1713260442
transform 1 0 1636 0 1 1305
box -2 -3 18 103
use MUX2X1  MUX2X1_19
timestamp 1713260442
transform 1 0 1652 0 1 1305
box -2 -3 50 103
use NAND2X1  NAND2X1_51
timestamp 1713260442
transform -1 0 1724 0 1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_59
timestamp 1713260442
transform -1 0 1756 0 1 1305
box -2 -3 34 103
use NAND3X1  NAND3X1_12
timestamp 1713260442
transform -1 0 1788 0 1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_62
timestamp 1713260442
transform 1 0 1788 0 1 1305
box -2 -3 26 103
use AND2X2  AND2X2_3
timestamp 1713260442
transform -1 0 1844 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_61
timestamp 1713260442
transform -1 0 1876 0 1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_66
timestamp 1713260442
transform -1 0 1900 0 1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_63
timestamp 1713260442
transform -1 0 1924 0 1 1305
box -2 -3 26 103
use NAND3X1  NAND3X1_13
timestamp 1713260442
transform -1 0 1956 0 1 1305
box -2 -3 34 103
use AOI21X1  AOI21X1_26
timestamp 1713260442
transform -1 0 1988 0 1 1305
box -2 -3 34 103
use XNOR2X1  XNOR2X1_7
timestamp 1713260442
transform -1 0 2044 0 1 1305
box -2 -3 58 103
use FILL  FILL_14_1
timestamp 1713260442
transform 1 0 2044 0 1 1305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_96
timestamp 1713260442
transform 1 0 4 0 -1 1505
box -2 -3 98 103
use OAI21X1  OAI21X1_40
timestamp 1713260442
transform 1 0 100 0 -1 1505
box -2 -3 34 103
use AOI21X1  AOI21X1_89
timestamp 1713260442
transform 1 0 132 0 -1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_43
timestamp 1713260442
transform 1 0 164 0 -1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_30
timestamp 1713260442
transform -1 0 220 0 -1 1505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_110
timestamp 1713260442
transform 1 0 220 0 -1 1505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_18
timestamp 1713260442
transform 1 0 316 0 -1 1505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_6
timestamp 1713260442
transform 1 0 412 0 -1 1505
box -2 -3 98 103
use FILL  FILL_14_0_0
timestamp 1713260442
transform -1 0 516 0 -1 1505
box -2 -3 10 103
use FILL  FILL_14_0_1
timestamp 1713260442
transform -1 0 524 0 -1 1505
box -2 -3 10 103
use INVX1  INVX1_40
timestamp 1713260442
transform -1 0 540 0 -1 1505
box -2 -3 18 103
use NAND2X1  NAND2X1_95
timestamp 1713260442
transform 1 0 540 0 -1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_163
timestamp 1713260442
transform -1 0 596 0 -1 1505
box -2 -3 34 103
use BUFX4  BUFX4_45
timestamp 1713260442
transform 1 0 596 0 -1 1505
box -2 -3 34 103
use INVX1  INVX1_22
timestamp 1713260442
transform 1 0 628 0 -1 1505
box -2 -3 18 103
use NOR2X1  NOR2X1_18
timestamp 1713260442
transform -1 0 668 0 -1 1505
box -2 -3 26 103
use DFFSR  DFFSR_4
timestamp 1713260442
transform -1 0 844 0 -1 1505
box -2 -3 178 103
use INVX1  INVX1_19
timestamp 1713260442
transform 1 0 844 0 -1 1505
box -2 -3 18 103
use OAI21X1  OAI21X1_162
timestamp 1713260442
transform 1 0 860 0 -1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_94
timestamp 1713260442
transform -1 0 916 0 -1 1505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_5
timestamp 1713260442
transform -1 0 1012 0 -1 1505
box -2 -3 98 103
use FILL  FILL_14_1_0
timestamp 1713260442
transform -1 0 1020 0 -1 1505
box -2 -3 10 103
use FILL  FILL_14_1_1
timestamp 1713260442
transform -1 0 1028 0 -1 1505
box -2 -3 10 103
use NAND3X1  NAND3X1_9
timestamp 1713260442
transform -1 0 1060 0 -1 1505
box -2 -3 34 103
use NAND3X1  NAND3X1_15
timestamp 1713260442
transform 1 0 1060 0 -1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_77
timestamp 1713260442
transform -1 0 1116 0 -1 1505
box -2 -3 26 103
use NAND2X1  NAND2X1_99
timestamp 1713260442
transform -1 0 1140 0 -1 1505
box -2 -3 26 103
use NAND3X1  NAND3X1_3
timestamp 1713260442
transform 1 0 1140 0 -1 1505
box -2 -3 34 103
use NAND3X1  NAND3X1_2
timestamp 1713260442
transform 1 0 1172 0 -1 1505
box -2 -3 34 103
use NAND3X1  NAND3X1_7
timestamp 1713260442
transform 1 0 1204 0 -1 1505
box -2 -3 34 103
use NAND3X1  NAND3X1_14
timestamp 1713260442
transform 1 0 1236 0 -1 1505
box -2 -3 34 103
use NAND3X1  NAND3X1_1
timestamp 1713260442
transform 1 0 1268 0 -1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_66
timestamp 1713260442
transform 1 0 1300 0 -1 1505
box -2 -3 26 103
use BUFX4  BUFX4_11
timestamp 1713260442
transform -1 0 1356 0 -1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_78
timestamp 1713260442
transform 1 0 1356 0 -1 1505
box -2 -3 26 103
use XNOR2X1  XNOR2X1_1
timestamp 1713260442
transform -1 0 1436 0 -1 1505
box -2 -3 58 103
use NAND2X1  NAND2X1_54
timestamp 1713260442
transform 1 0 1436 0 -1 1505
box -2 -3 26 103
use NAND2X1  NAND2X1_61
timestamp 1713260442
transform 1 0 1460 0 -1 1505
box -2 -3 26 103
use AOI21X1  AOI21X1_25
timestamp 1713260442
transform 1 0 1484 0 -1 1505
box -2 -3 34 103
use FILL  FILL_14_2_0
timestamp 1713260442
transform -1 0 1524 0 -1 1505
box -2 -3 10 103
use FILL  FILL_14_2_1
timestamp 1713260442
transform -1 0 1532 0 -1 1505
box -2 -3 10 103
use AOI22X1  AOI22X1_1
timestamp 1713260442
transform -1 0 1572 0 -1 1505
box -2 -3 42 103
use OAI21X1  OAI21X1_58
timestamp 1713260442
transform -1 0 1604 0 -1 1505
box -2 -3 34 103
use INVX1  INVX1_9
timestamp 1713260442
transform 1 0 1604 0 -1 1505
box -2 -3 18 103
use NAND2X1  NAND2X1_64
timestamp 1713260442
transform 1 0 1620 0 -1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_60
timestamp 1713260442
transform 1 0 1644 0 -1 1505
box -2 -3 34 103
use AOI22X1  AOI22X1_2
timestamp 1713260442
transform -1 0 1716 0 -1 1505
box -2 -3 42 103
use NAND2X1  NAND2X1_55
timestamp 1713260442
transform 1 0 1716 0 -1 1505
box -2 -3 26 103
use AOI21X1  AOI21X1_27
timestamp 1713260442
transform -1 0 1772 0 -1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_65
timestamp 1713260442
transform 1 0 1772 0 -1 1505
box -2 -3 26 103
use NOR2X1  NOR2X1_26
timestamp 1713260442
transform -1 0 1820 0 -1 1505
box -2 -3 26 103
use AOI22X1  AOI22X1_3
timestamp 1713260442
transform 1 0 1820 0 -1 1505
box -2 -3 42 103
use NOR2X1  NOR2X1_36
timestamp 1713260442
transform -1 0 1884 0 -1 1505
box -2 -3 26 103
use NAND2X1  NAND2X1_53
timestamp 1713260442
transform 1 0 1884 0 -1 1505
box -2 -3 26 103
use NOR2X1  NOR2X1_27
timestamp 1713260442
transform 1 0 1908 0 -1 1505
box -2 -3 26 103
use NAND3X1  NAND3X1_6
timestamp 1713260442
transform 1 0 1932 0 -1 1505
box -2 -3 34 103
use NAND3X1  NAND3X1_5
timestamp 1713260442
transform -1 0 1996 0 -1 1505
box -2 -3 34 103
use AND2X2  AND2X2_2
timestamp 1713260442
transform -1 0 2028 0 -1 1505
box -2 -3 34 103
use BUFX2  BUFX2_11
timestamp 1713260442
transform -1 0 2052 0 -1 1505
box -2 -3 26 103
use BUFX2  BUFX2_2
timestamp 1713260442
transform -1 0 28 0 1 1505
box -2 -3 26 103
use BUFX2  BUFX2_1
timestamp 1713260442
transform -1 0 52 0 1 1505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_22
timestamp 1713260442
transform 1 0 52 0 1 1505
box -2 -3 98 103
use NOR2X1  NOR2X1_63
timestamp 1713260442
transform 1 0 148 0 1 1505
box -2 -3 26 103
use DFFSR  DFFSR_9
timestamp 1713260442
transform -1 0 348 0 1 1505
box -2 -3 178 103
use DFFSR  DFFSR_15
timestamp 1713260442
transform -1 0 180 0 -1 1705
box -2 -3 178 103
use DFFSR  DFFSR_13
timestamp 1713260442
transform -1 0 356 0 -1 1705
box -2 -3 178 103
use AOI21X1  AOI21X1_86
timestamp 1713260442
transform 1 0 348 0 1 1505
box -2 -3 34 103
use DFFSR  DFFSR_12
timestamp 1713260442
transform -1 0 532 0 -1 1705
box -2 -3 178 103
use NOR2X1  NOR2X1_60
timestamp 1713260442
transform -1 0 404 0 1 1505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_38
timestamp 1713260442
transform 1 0 404 0 1 1505
box -2 -3 98 103
use FILL  FILL_15_0_0
timestamp 1713260442
transform 1 0 500 0 1 1505
box -2 -3 10 103
use FILL  FILL_15_0_1
timestamp 1713260442
transform 1 0 508 0 1 1505
box -2 -3 10 103
use OAI21X1  OAI21X1_6
timestamp 1713260442
transform 1 0 516 0 1 1505
box -2 -3 34 103
use FILL  FILL_16_0_0
timestamp 1713260442
transform -1 0 540 0 -1 1705
box -2 -3 10 103
use FILL  FILL_16_0_1
timestamp 1713260442
transform -1 0 548 0 -1 1705
box -2 -3 10 103
use AOI21X1  AOI21X1_14
timestamp 1713260442
transform 1 0 636 0 -1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_37
timestamp 1713260442
transform -1 0 636 0 -1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_34
timestamp 1713260442
transform 1 0 580 0 -1 1705
box -2 -3 34 103
use BUFX4  BUFX4_14
timestamp 1713260442
transform -1 0 580 0 -1 1705
box -2 -3 34 103
use AOI21X1  AOI21X1_15
timestamp 1713260442
transform 1 0 572 0 1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_6
timestamp 1713260442
transform 1 0 548 0 1 1505
box -2 -3 26 103
use NOR2X1  NOR2X1_17
timestamp 1713260442
transform -1 0 692 0 -1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_39
timestamp 1713260442
transform 1 0 700 0 1 1505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_95
timestamp 1713260442
transform 1 0 692 0 -1 1705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_46
timestamp 1713260442
transform 1 0 604 0 1 1505
box -2 -3 98 103
use NAND2X1  NAND2X1_42
timestamp 1713260442
transform -1 0 756 0 1 1505
box -2 -3 26 103
use NAND2X1  NAND2X1_59
timestamp 1713260442
transform 1 0 756 0 1 1505
box -2 -3 26 103
use DFFSR  DFFSR_8
timestamp 1713260442
transform 1 0 780 0 1 1505
box -2 -3 178 103
use OAI21X1  OAI21X1_2
timestamp 1713260442
transform 1 0 788 0 -1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_2
timestamp 1713260442
transform -1 0 844 0 -1 1705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_34
timestamp 1713260442
transform -1 0 940 0 -1 1705
box -2 -3 98 103
use XNOR2X1  XNOR2X1_4
timestamp 1713260442
transform 1 0 940 0 -1 1705
box -2 -3 58 103
use OAI21X1  OAI21X1_55
timestamp 1713260442
transform -1 0 988 0 1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_28
timestamp 1713260442
transform -1 0 1052 0 -1 1705
box -2 -3 26 103
use FILL  FILL_16_1_1
timestamp 1713260442
transform -1 0 1028 0 -1 1705
box -2 -3 10 103
use FILL  FILL_16_1_0
timestamp 1713260442
transform -1 0 1020 0 -1 1705
box -2 -3 10 103
use INVX2  INVX2_2
timestamp 1713260442
transform -1 0 1012 0 -1 1705
box -2 -3 18 103
use INVX1  INVX1_3
timestamp 1713260442
transform 1 0 1028 0 1 1505
box -2 -3 18 103
use FILL  FILL_15_1_1
timestamp 1713260442
transform 1 0 1020 0 1 1505
box -2 -3 10 103
use FILL  FILL_15_1_0
timestamp 1713260442
transform 1 0 1012 0 1 1505
box -2 -3 10 103
use NOR2X1  NOR2X1_34
timestamp 1713260442
transform -1 0 1012 0 1 1505
box -2 -3 26 103
use NOR2X1  NOR2X1_2
timestamp 1713260442
transform -1 0 1100 0 -1 1705
box -2 -3 26 103
use NAND2X1  NAND2X1_58
timestamp 1713260442
transform 1 0 1052 0 -1 1705
box -2 -3 26 103
use NAND2X1  NAND2X1_88
timestamp 1713260442
transform 1 0 1068 0 1 1505
box -2 -3 26 103
use NOR2X1  NOR2X1_56
timestamp 1713260442
transform 1 0 1044 0 1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_53
timestamp 1713260442
transform 1 0 1180 0 -1 1705
box -2 -3 34 103
use NAND3X1  NAND3X1_4
timestamp 1713260442
transform 1 0 1148 0 -1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_10
timestamp 1713260442
transform -1 0 1148 0 -1 1705
box -2 -3 26 103
use NOR2X1  NOR2X1_12
timestamp 1713260442
transform -1 0 1124 0 -1 1705
box -2 -3 26 103
use NOR2X1  NOR2X1_21
timestamp 1713260442
transform 1 0 1172 0 1 1505
box -2 -3 26 103
use NAND2X1  NAND2X1_11
timestamp 1713260442
transform 1 0 1148 0 1 1505
box -2 -3 26 103
use BUFX4  BUFX4_15
timestamp 1713260442
transform 1 0 1116 0 1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_58
timestamp 1713260442
transform 1 0 1092 0 1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_54
timestamp 1713260442
transform -1 0 1292 0 -1 1705
box -2 -3 34 103
use NOR2X1  NOR2X1_32
timestamp 1713260442
transform 1 0 1236 0 -1 1705
box -2 -3 26 103
use NOR2X1  NOR2X1_57
timestamp 1713260442
transform 1 0 1212 0 -1 1705
box -2 -3 26 103
use NAND2X1  NAND2X1_100
timestamp 1713260442
transform 1 0 1220 0 1 1505
box -2 -3 26 103
use NAND2X1  NAND2X1_89
timestamp 1713260442
transform 1 0 1196 0 1 1505
box -2 -3 26 103
use DFFSR  DFFSR_1
timestamp 1713260442
transform -1 0 1420 0 1 1505
box -2 -3 178 103
use DFFSR  DFFSR_19
timestamp 1713260442
transform -1 0 1596 0 1 1505
box -2 -3 178 103
use XNOR2X1  XNOR2X1_3
timestamp 1713260442
transform 1 0 1292 0 -1 1705
box -2 -3 58 103
use DFFSR  DFFSR_5
timestamp 1713260442
transform -1 0 1524 0 -1 1705
box -2 -3 178 103
use FILL  FILL_15_2_0
timestamp 1713260442
transform 1 0 1596 0 1 1505
box -2 -3 10 103
use FILL  FILL_15_2_1
timestamp 1713260442
transform 1 0 1604 0 1 1505
box -2 -3 10 103
use DFFSR  DFFSR_21
timestamp 1713260442
transform 1 0 1612 0 1 1505
box -2 -3 178 103
use FILL  FILL_16_2_0
timestamp 1713260442
transform -1 0 1532 0 -1 1705
box -2 -3 10 103
use FILL  FILL_16_2_1
timestamp 1713260442
transform -1 0 1540 0 -1 1705
box -2 -3 10 103
use XNOR2X1  XNOR2X1_6
timestamp 1713260442
transform -1 0 1596 0 -1 1705
box -2 -3 58 103
use XNOR2X1  XNOR2X1_5
timestamp 1713260442
transform 1 0 1596 0 -1 1705
box -2 -3 58 103
use NOR2X1  NOR2X1_35
timestamp 1713260442
transform -1 0 1812 0 1 1505
box -2 -3 26 103
use NOR2X1  NOR2X1_37
timestamp 1713260442
transform -1 0 1836 0 1 1505
box -2 -3 26 103
use DFFSR  DFFSR_20
timestamp 1713260442
transform 1 0 1652 0 -1 1705
box -2 -3 178 103
use AOI21X1  AOI21X1_24
timestamp 1713260442
transform 1 0 1884 0 -1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_57
timestamp 1713260442
transform -1 0 1884 0 -1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_60
timestamp 1713260442
transform 1 0 1828 0 -1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_49
timestamp 1713260442
transform 1 0 1884 0 1 1505
box -2 -3 34 103
use INVX1  INVX1_8
timestamp 1713260442
transform 1 0 1868 0 1 1505
box -2 -3 18 103
use OAI21X1  OAI21X1_50
timestamp 1713260442
transform 1 0 1836 0 1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_56
timestamp 1713260442
transform 1 0 1972 0 -1 1705
box -2 -3 34 103
use XOR2X1  XOR2X1_1
timestamp 1713260442
transform 1 0 1916 0 -1 1705
box -2 -3 58 103
use AND2X2  AND2X2_1
timestamp 1713260442
transform -1 0 1948 0 1 1505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_70
timestamp 1713260442
transform 1 0 1948 0 1 1505
box -2 -3 98 103
use FILL  FILL_16_1
timestamp 1713260442
transform 1 0 2044 0 1 1505
box -2 -3 10 103
use NAND3X1  NAND3X1_11
timestamp 1713260442
transform 1 0 2004 0 -1 1705
box -2 -3 34 103
use INVX1  INVX1_7
timestamp 1713260442
transform -1 0 2052 0 -1 1705
box -2 -3 18 103
use BUFX2  BUFX2_7
timestamp 1713260442
transform -1 0 28 0 1 1705
box -2 -3 26 103
use BUFX2  BUFX2_8
timestamp 1713260442
transform -1 0 52 0 1 1705
box -2 -3 26 103
use CLKBUF1  CLKBUF1_8
timestamp 1713260442
transform 1 0 52 0 1 1705
box -2 -3 74 103
use BUFX2  BUFX2_5
timestamp 1713260442
transform -1 0 148 0 1 1705
box -2 -3 26 103
use BUFX2  BUFX2_4
timestamp 1713260442
transform -1 0 172 0 1 1705
box -2 -3 26 103
use BUFX2  BUFX2_6
timestamp 1713260442
transform -1 0 196 0 1 1705
box -2 -3 26 103
use DFFSR  DFFSR_14
timestamp 1713260442
transform -1 0 372 0 1 1705
box -2 -3 178 103
use BUFX4  BUFX4_12
timestamp 1713260442
transform -1 0 404 0 1 1705
box -2 -3 34 103
use BUFX2  BUFX2_3
timestamp 1713260442
transform -1 0 428 0 1 1705
box -2 -3 26 103
use FILL  FILL_17_0_0
timestamp 1713260442
transform -1 0 436 0 1 1705
box -2 -3 10 103
use FILL  FILL_17_0_1
timestamp 1713260442
transform -1 0 444 0 1 1705
box -2 -3 10 103
use DFFSR  DFFSR_11
timestamp 1713260442
transform -1 0 620 0 1 1705
box -2 -3 178 103
use DFFPOSX1  DFFPOSX1_90
timestamp 1713260442
transform -1 0 716 0 1 1705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_45
timestamp 1713260442
transform -1 0 812 0 1 1705
box -2 -3 98 103
use INVX8  INVX8_1
timestamp 1713260442
transform 1 0 812 0 1 1705
box -2 -3 42 103
use CLKBUF1  CLKBUF1_6
timestamp 1713260442
transform -1 0 924 0 1 1705
box -2 -3 74 103
use DFFSR  DFFSR_7
timestamp 1713260442
transform 1 0 924 0 1 1705
box -2 -3 178 103
use FILL  FILL_17_1_0
timestamp 1713260442
transform 1 0 1100 0 1 1705
box -2 -3 10 103
use FILL  FILL_17_1_1
timestamp 1713260442
transform 1 0 1108 0 1 1705
box -2 -3 10 103
use BUFX4  BUFX4_13
timestamp 1713260442
transform 1 0 1116 0 1 1705
box -2 -3 34 103
use CLKBUF1  CLKBUF1_3
timestamp 1713260442
transform -1 0 1220 0 1 1705
box -2 -3 74 103
use NOR2X1  NOR2X1_33
timestamp 1713260442
transform 1 0 1220 0 1 1705
box -2 -3 26 103
use INVX1  INVX1_4
timestamp 1713260442
transform -1 0 1260 0 1 1705
box -2 -3 18 103
use NOR2X1  NOR2X1_29
timestamp 1713260442
transform -1 0 1284 0 1 1705
box -2 -3 26 103
use INVX2  INVX2_3
timestamp 1713260442
transform -1 0 1300 0 1 1705
box -2 -3 18 103
use DFFSR  DFFSR_6
timestamp 1713260442
transform -1 0 1476 0 1 1705
box -2 -3 178 103
use FILL  FILL_17_2_0
timestamp 1713260442
transform 1 0 1476 0 1 1705
box -2 -3 10 103
use FILL  FILL_17_2_1
timestamp 1713260442
transform 1 0 1484 0 1 1705
box -2 -3 10 103
use DFFSR  DFFSR_17
timestamp 1713260442
transform 1 0 1492 0 1 1705
box -2 -3 178 103
use CLKBUF1  CLKBUF1_2
timestamp 1713260442
transform 1 0 1668 0 1 1705
box -2 -3 74 103
use DFFSR  DFFSR_18
timestamp 1713260442
transform 1 0 1740 0 1 1705
box -2 -3 178 103
use INVX1  INVX1_6
timestamp 1713260442
transform -1 0 1932 0 1 1705
box -2 -3 18 103
use NAND3X1  NAND3X1_10
timestamp 1713260442
transform 1 0 1932 0 1 1705
box -2 -3 34 103
use INVX1  INVX1_1
timestamp 1713260442
transform 1 0 1964 0 1 1705
box -2 -3 18 103
use BUFX2  BUFX2_15
timestamp 1713260442
transform 1 0 1980 0 1 1705
box -2 -3 26 103
use INVX1  INVX1_2
timestamp 1713260442
transform 1 0 2004 0 1 1705
box -2 -3 18 103
use BUFX2  BUFX2_9
timestamp 1713260442
transform 1 0 2020 0 1 1705
box -2 -3 26 103
use FILL  FILL_18_1
timestamp 1713260442
transform 1 0 2044 0 1 1705
box -2 -3 10 103
<< labels >>
flabel metal6 s 496 -30 512 -22 7 FreeSans 24 270 0 0 vdd
port 0 nsew
flabel metal6 s 1016 -30 1032 -22 7 FreeSans 24 270 0 0 gnd
port 1 nsew
flabel metal2 s 118 1828 122 1832 3 FreeSans 24 90 0 0 clk
port 2 nsew
flabel metal2 s 830 1828 834 1832 3 FreeSans 24 90 0 0 reset
port 3 nsew
flabel metal3 s 2078 58 2082 62 3 FreeSans 24 270 0 0 d_in[0]
port 4 nsew
flabel metal3 s 2078 448 2082 452 3 FreeSans 24 0 0 0 d_in[1]
port 5 nsew
flabel metal3 s 2078 468 2082 472 3 FreeSans 24 0 0 0 d_in[2]
port 6 nsew
flabel metal3 s 2078 548 2082 552 3 FreeSans 24 0 0 0 d_in[3]
port 7 nsew
flabel metal3 s 2078 1048 2082 1052 3 FreeSans 24 0 0 0 d_in[4]
port 8 nsew
flabel metal3 s 2078 1248 2082 1252 3 FreeSans 24 0 0 0 d_in[5]
port 9 nsew
flabel metal3 s 2078 1268 2082 1272 3 FreeSans 24 0 0 0 d_in[6]
port 10 nsew
flabel metal3 s 2078 1308 2082 1312 3 FreeSans 24 0 0 0 d_in[7]
port 11 nsew
flabel metal2 s 1934 1828 1938 1832 3 FreeSans 24 90 0 0 wr_en
port 12 nsew
flabel metal2 s 1958 1828 1962 1832 3 FreeSans 24 90 0 0 rd_en
port 13 nsew
flabel metal3 s 2078 1768 2082 1772 3 FreeSans 24 90 0 0 full
port 14 nsew
flabel metal3 s 2078 1748 2082 1752 3 FreeSans 24 90 0 0 empty
port 15 nsew
flabel metal3 s -26 1548 -22 1552 7 FreeSans 24 0 0 0 d_out[0]
port 16 nsew
flabel metal3 s -26 1568 -22 1572 7 FreeSans 24 0 0 0 d_out[1]
port 17 nsew
flabel metal3 s -26 1718 -22 1722 7 FreeSans 24 0 0 0 d_out[2]
port 18 nsew
flabel metal3 s -26 1738 -22 1742 7 FreeSans 24 90 0 0 d_out[3]
port 19 nsew
flabel metal3 s -26 1758 -22 1762 7 FreeSans 24 90 0 0 d_out[4]
port 20 nsew
flabel metal3 s -26 1778 -22 1782 7 FreeSans 24 90 0 0 d_out[5]
port 21 nsew
flabel metal3 s -26 1798 -22 1802 7 FreeSans 24 90 0 0 d_out[6]
port 22 nsew
flabel metal3 s -26 1818 -22 1822 7 FreeSans 24 90 0 0 d_out[7]
port 23 nsew
flabel metal2 s 1990 -22 1994 -18 3 FreeSans 24 270 0 0 fifo_counter[0]
port 24 nsew
flabel metal2 s 2014 -22 2018 -18 3 FreeSans 24 270 0 0 fifo_counter[1]
port 25 nsew
flabel metal2 s 2030 -22 2034 -18 3 FreeSans 24 270 0 0 fifo_counter[2]
port 26 nsew
flabel metal2 s 2046 -22 2050 -18 3 FreeSans 24 270 0 0 fifo_counter[3]
port 27 nsew
flabel metal2 s 2062 -22 2066 -18 3 FreeSans 24 270 0 0 fifo_counter[4]
port 28 nsew
<< end >>
